// Benchmark "i10" written by ABC on Fri Mar 11 15:18:06 2022

module i10 ( 
    \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) , \V10(0) ,
    \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) , \V248(0) ,
    \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) , \V66(0) ,
    \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) , \V45(0) ,
    \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) , \V34(0) ,
    \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) , \V293(0) ,
    \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) , \V275(0) ,
    \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) , \V257(4) ,
    \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) , \V149(3) ,
    \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) , \V165(6) ,
    \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) , \V169(0) ,
    \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) , \V165(3) ,
    \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) , \V288(4) ,
    \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) , \V229(3) ,
    \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) , \V223(3) ,
    \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) , \V189(3) ,
    \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) , \V183(3) ,
    \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) , \V239(2) ,
    \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) , \V234(1) ,
    \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) , \V199(0) ,
    \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) , \V257(0) ,
    \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) , \V32(10) ,
    \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) , \V84(2) ,
    \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) , \V14(0) ,
    \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) , \V213(1) ,
    \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) , \V8(0) ,
    \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) ,
    \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) ,
    \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) ,
    \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) ,
    \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) ,
    \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) ,
    \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) ,
    \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) ,
    \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) ,
    \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) ,
    \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) ,
    \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) ,
    \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) ,
    \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) ,
    \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) ,
    \V78(0) , \V94(0) , \V94(1) ,
    \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) ,
    \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) ,
    V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546,
    V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) ,
    \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587,
    \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630,
    \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781,
    V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) ,
    \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) ,
    \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) ,
    \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) ,
    \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) ,
    \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) ,
    \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378,
    V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) ,
    \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) ,
    \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539,
    \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) ,
    \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) ,
    \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) ,
    V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) ,
    \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) ,
    \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) ,
    \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832,
    \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) ,
    \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) ,
    \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) ,
    \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) ,
    \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653,
    V654, V655, V656, V1370, V1371, V1372, V1373, V1374  );
  input  \V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) ,
    \V10(0) , \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) ,
    \V248(0) , \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) ,
    \V66(0) , \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) ,
    \V45(0) , \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) ,
    \V34(0) , \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) ,
    \V293(0) , \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) ,
    \V275(0) , \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) ,
    \V257(4) , \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) ,
    \V149(3) , \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) ,
    \V165(6) , \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) ,
    \V169(0) , \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) ,
    \V165(3) , \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) ,
    \V288(4) , \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) ,
    \V229(3) , \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) ,
    \V223(3) , \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) ,
    \V189(3) , \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) ,
    \V183(3) , \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) ,
    \V239(2) , \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) ,
    \V234(1) , \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) ,
    \V199(0) , \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) ,
    \V257(0) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) ,
    \V32(10) , \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) ,
    \V84(2) , \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) ,
    \V14(0) , \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) ,
    \V213(1) , \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) ,
    \V8(0) , \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) ,
    \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) ,
    \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) ,
    \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) ,
    \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) ,
    \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) ,
    \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) ,
    \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) ,
    \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) ,
    \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) ,
    \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) ,
    \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) ,
    \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) ,
    \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) ,
    \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) ,
    \V78(0) , \V94(0) , \V94(1) ;
  output \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) ,
    \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) ,
    V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546,
    V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) ,
    \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587,
    \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630,
    \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781,
    V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) ,
    \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) ,
    \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) ,
    \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) ,
    \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) ,
    \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263,
    V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) ,
    \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378,
    V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428,
    V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) ,
    \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) ,
    \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539,
    \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) ,
    \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) ,
    \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) ,
    V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) ,
    \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) ,
    \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) ,
    \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832,
    \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) ,
    \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) ,
    \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) ,
    \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) ,
    \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653,
    V654, V655, V656, V1370, V1371, V1372, V1373, V1374;
  wire new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n904_,
    new_n905_, new_n906_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1096_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1109_, new_n1110_,
    new_n1112_, new_n1113_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1123_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1371_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1378_,
    new_n1379_, new_n1380_, new_n1382_, new_n1383_, new_n1384_, new_n1386_,
    new_n1387_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1395_, new_n1396_, new_n1398_, new_n1399_, new_n1401_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1435_, new_n1436_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1443_, new_n1447_,
    new_n1448_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1497_, new_n1498_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1523_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1565_, new_n1567_, new_n1569_,
    new_n1571_, new_n1573_, new_n1575_, new_n1576_, new_n1579_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1589_, new_n1590_, new_n1591_, new_n1593_, new_n1595_, new_n1597_,
    new_n1598_, new_n1599_, new_n1601_, new_n1607_, new_n1608_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1634_, new_n1635_, new_n1637_, new_n1638_, new_n1639_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1654_, new_n1655_,
    new_n1656_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1665_, new_n1666_, new_n1667_, new_n1669_, new_n1671_,
    new_n1673_, new_n1674_, new_n1675_, new_n1677_, new_n1678_, new_n1679_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1751_, new_n1752_, new_n1754_, new_n1755_, new_n1757_, new_n1758_,
    new_n1759_, new_n1761_, new_n1762_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1769_, new_n1770_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1779_, new_n1780_, new_n1782_,
    new_n1783_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1791_, new_n1792_, new_n1794_, new_n1795_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1822_, new_n1824_, new_n1826_, new_n1828_, new_n1830_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1837_, new_n1838_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1850_, new_n1852_,
    new_n1853_, new_n1855_, new_n1857_, new_n1858_, new_n1862_, new_n1864_,
    new_n1866_, new_n1868_, new_n1870_, new_n1872_, new_n1875_, new_n1876_,
    new_n1879_, new_n1880_, new_n1881_, new_n1884_, new_n1887_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1907_, new_n1908_, new_n1909_, new_n1911_,
    new_n1912_, new_n1914_, new_n1915_, new_n1917_, new_n1919_, new_n1921_,
    new_n1923_, new_n1927_, new_n1929_, new_n1931_;
  INVX1    g0000(.A(\V53(0) ), .Y(new_n482_));
  INVX1    g0001(.A(\V149(1) ), .Y(new_n483_));
  INVX1    g0002(.A(\V149(2) ), .Y(new_n484_));
  INVX1    g0003(.A(\V149(3) ), .Y(new_n485_));
  NOR4X1   g0004(.A(new_n485_), .B(new_n484_), .C(new_n483_), .D(\V149(0) ), .Y(new_n486_));
  INVX1    g0005(.A(\V169(0) ), .Y(new_n487_));
  INVX1    g0006(.A(\V165(6) ), .Y(new_n488_));
  INVX1    g0007(.A(\V70(0) ), .Y(new_n489_));
  INVX1    g0008(.A(\V165(3) ), .Y(new_n490_));
  NOR4X1   g0009(.A(new_n490_), .B(\V165(5) ), .C(\V165(4) ), .D(new_n489_), .Y(new_n491_));
  AND2X1   g0010(.A(new_n491_), .B(new_n488_), .Y(new_n492_));
  NOR2X1   g0011(.A(\V51(0) ), .B(\V52(0) ), .Y(new_n493_));
  INVX1    g0012(.A(new_n493_), .Y(\V802(0) ));
  INVX1    g0013(.A(\V149(6) ), .Y(new_n495_));
  INVX1    g0014(.A(\V149(4) ), .Y(new_n496_));
  INVX1    g0015(.A(\V149(0) ), .Y(new_n497_));
  NAND3X1  g0016(.A(new_n484_), .B(\V149(1) ), .C(new_n497_), .Y(new_n498_));
  NAND3X1  g0017(.A(new_n485_), .B(\V149(5) ), .C(\V149(7) ), .Y(new_n499_));
  OR4X1    g0018(.A(new_n499_), .B(new_n498_), .C(new_n496_), .D(new_n495_), .Y(new_n500_));
  INVX1    g0019(.A(\V149(7) ), .Y(new_n501_));
  NAND3X1  g0020(.A(new_n485_), .B(\V149(5) ), .C(new_n501_), .Y(new_n502_));
  OR4X1    g0021(.A(new_n502_), .B(new_n498_), .C(new_n496_), .D(new_n495_), .Y(new_n503_));
  AND2X1   g0022(.A(new_n503_), .B(new_n500_), .Y(new_n504_));
  NOR3X1   g0023(.A(new_n504_), .B(\V802(0) ), .C(\V55(0) ), .Y(new_n505_));
  OR4X1    g0024(.A(new_n484_), .B(new_n483_), .C(\V149(0) ), .D(new_n496_), .Y(new_n506_));
  NOR2X1   g0025(.A(new_n506_), .B(\V149(3) ), .Y(new_n507_));
  NOR3X1   g0026(.A(\V149(2) ), .B(\V149(1) ), .C(\V149(0) ), .Y(new_n508_));
  NOR3X1   g0027(.A(new_n508_), .B(new_n507_), .C(new_n505_), .Y(new_n509_));
  OR4X1    g0028(.A(new_n509_), .B(new_n492_), .C(\V291(0) ), .D(new_n487_), .Y(new_n510_));
  INVX1    g0029(.A(\V165(0) ), .Y(new_n511_));
  INVX1    g0030(.A(\V165(2) ), .Y(new_n512_));
  INVX1    g0031(.A(\V165(1) ), .Y(new_n513_));
  INVX1    g0032(.A(\V165(4) ), .Y(new_n514_));
  NAND4X1  g0033(.A(\V261(0) ), .B(\V165(7) ), .C(\V165(5) ), .D(\V70(0) ), .Y(new_n515_));
  OR4X1    g0034(.A(new_n515_), .B(new_n490_), .C(new_n488_), .D(new_n514_), .Y(new_n516_));
  OR4X1    g0035(.A(new_n516_), .B(new_n513_), .C(new_n512_), .D(new_n511_), .Y(new_n517_));
  NOR3X1   g0036(.A(new_n517_), .B(new_n510_), .C(\V292(0) ), .Y(new_n518_));
  INVX1    g0037(.A(\V261(0) ), .Y(\V1833(0) ));
  NAND4X1  g0038(.A(\V165(3) ), .B(\V165(7) ), .C(\V165(6) ), .D(\V165(5) ), .Y(new_n520_));
  OR4X1    g0039(.A(new_n520_), .B(\V1833(0) ), .C(\V204(0) ), .D(new_n514_), .Y(new_n521_));
  NOR4X1   g0040(.A(new_n521_), .B(new_n513_), .C(new_n512_), .D(new_n511_), .Y(new_n522_));
  OR2X1    g0041(.A(\V149(0) ), .B(\V149(4) ), .Y(new_n523_));
  NOR4X1   g0042(.A(new_n523_), .B(\V149(3) ), .C(new_n484_), .D(new_n483_), .Y(new_n524_));
  OR4X1    g0043(.A(new_n524_), .B(new_n522_), .C(new_n518_), .D(\V262(0) ), .Y(new_n525_));
  OR4X1    g0044(.A(new_n525_), .B(new_n486_), .C(new_n482_), .D(\V56(0) ), .Y(new_n526_));
  INVX1    g0045(.A(\V149(5) ), .Y(new_n527_));
  NAND3X1  g0046(.A(new_n485_), .B(new_n527_), .C(\V149(7) ), .Y(new_n528_));
  NOR4X1   g0047(.A(new_n528_), .B(new_n498_), .C(new_n496_), .D(new_n495_), .Y(new_n529_));
  INVX1    g0048(.A(new_n529_), .Y(new_n530_));
  INVX1    g0049(.A(\V56(0) ), .Y(new_n531_));
  INVX1    g0050(.A(\V57(0) ), .Y(new_n532_));
  NAND3X1  g0051(.A(new_n532_), .B(new_n482_), .C(new_n531_), .Y(new_n533_));
  INVX1    g0052(.A(\V169(1) ), .Y(new_n534_));
  OR2X1    g0053(.A(\V149(1) ), .B(\V149(0) ), .Y(new_n535_));
  OR4X1    g0054(.A(\V149(2) ), .B(\V149(1) ), .C(\V149(0) ), .D(\V174(0) ), .Y(new_n536_));
  NOR4X1   g0055(.A(new_n536_), .B(new_n535_), .C(new_n534_), .D(new_n485_), .Y(new_n537_));
  NOR2X1   g0056(.A(new_n535_), .B(new_n534_), .Y(new_n538_));
  INVX1    g0057(.A(new_n538_), .Y(new_n539_));
  INVX1    g0058(.A(\V88(2) ), .Y(new_n540_));
  OR2X1    g0059(.A(new_n536_), .B(\V149(3) ), .Y(new_n541_));
  OR4X1    g0060(.A(new_n541_), .B(new_n540_), .C(\V149(4) ), .D(\V149(5) ), .Y(new_n542_));
  OR4X1    g0061(.A(new_n536_), .B(\V149(3) ), .C(new_n496_), .D(new_n527_), .Y(new_n543_));
  OAI21X1  g0062(.A0(new_n542_), .A1(\V88(3) ), .B0(new_n543_), .Y(new_n544_));
  OR4X1    g0063(.A(new_n536_), .B(\V149(3) ), .C(\V149(4) ), .D(new_n527_), .Y(new_n545_));
  OR2X1    g0064(.A(new_n545_), .B(new_n540_), .Y(new_n546_));
  OR2X1    g0065(.A(new_n545_), .B(\V88(2) ), .Y(new_n547_));
  AOI21X1  g0066(.A0(new_n547_), .A1(new_n546_), .B0(\V88(3) ), .Y(new_n548_));
  INVX1    g0067(.A(\V88(3) ), .Y(new_n549_));
  AOI21X1  g0068(.A0(new_n547_), .A1(new_n542_), .B0(new_n549_), .Y(new_n550_));
  OR4X1    g0069(.A(new_n536_), .B(\V149(3) ), .C(new_n496_), .D(\V149(5) ), .Y(new_n551_));
  OR4X1    g0070(.A(new_n541_), .B(\V88(2) ), .C(\V149(4) ), .D(\V149(5) ), .Y(new_n552_));
  OAI21X1  g0071(.A0(new_n552_), .A1(new_n549_), .B0(new_n551_), .Y(new_n553_));
  NOR4X1   g0072(.A(new_n553_), .B(new_n550_), .C(new_n548_), .D(new_n544_), .Y(new_n554_));
  NOR2X1   g0073(.A(new_n554_), .B(new_n539_), .Y(new_n555_));
  OAI22X1  g0074(.A0(new_n555_), .A1(new_n537_), .B0(\V60(0) ), .B1(\V56(0) ), .Y(new_n556_));
  NOR2X1   g0075(.A(new_n536_), .B(new_n485_), .Y(new_n557_));
  INVX1    g0076(.A(new_n557_), .Y(new_n558_));
  OR4X1    g0077(.A(new_n485_), .B(new_n484_), .C(\V149(1) ), .D(\V149(0) ), .Y(new_n559_));
  AND2X1   g0078(.A(new_n559_), .B(new_n554_), .Y(new_n560_));
  INVX1    g0079(.A(\V278(0) ), .Y(new_n561_));
  NOR3X1   g0080(.A(new_n506_), .B(\V149(3) ), .C(\V174(0) ), .Y(new_n562_));
  OAI21X1  g0081(.A0(new_n561_), .A1(\V277(0) ), .B0(new_n562_), .Y(new_n563_));
  NAND3X1  g0082(.A(\V149(2) ), .B(new_n483_), .C(new_n497_), .Y(new_n564_));
  NOR3X1   g0083(.A(new_n564_), .B(\V149(3) ), .C(new_n527_), .Y(new_n565_));
  NOR3X1   g0084(.A(new_n564_), .B(\V149(3) ), .C(\V149(5) ), .Y(new_n566_));
  AOI21X1  g0085(.A0(new_n565_), .A1(new_n496_), .B0(new_n566_), .Y(new_n567_));
  NAND4X1  g0086(.A(new_n567_), .B(new_n563_), .C(new_n560_), .D(new_n558_), .Y(new_n568_));
  NAND3X1  g0087(.A(new_n568_), .B(new_n556_), .C(new_n533_), .Y(new_n569_));
  AND2X1   g0088(.A(new_n569_), .B(new_n530_), .Y(new_n570_));
  AND2X1   g0089(.A(new_n570_), .B(new_n526_), .Y(new_n571_));
  OR2X1    g0090(.A(new_n510_), .B(\V292(0) ), .Y(new_n572_));
  INVX1    g0091(.A(new_n517_), .Y(new_n573_));
  NOR4X1   g0092(.A(new_n522_), .B(new_n573_), .C(new_n572_), .D(\V262(0) ), .Y(new_n574_));
  INVX1    g0093(.A(new_n574_), .Y(new_n575_));
  INVX1    g0094(.A(\V262(0) ), .Y(new_n576_));
  NOR2X1   g0095(.A(new_n522_), .B(new_n518_), .Y(new_n577_));
  NAND2X1  g0096(.A(new_n577_), .B(new_n576_), .Y(new_n578_));
  INVX1    g0097(.A(new_n486_), .Y(new_n579_));
  AOI21X1  g0098(.A0(new_n562_), .A1(\V277(0) ), .B0(new_n561_), .Y(new_n580_));
  NOR2X1   g0099(.A(\V60(0) ), .B(\V59(0) ), .Y(new_n581_));
  NOR3X1   g0100(.A(new_n581_), .B(new_n580_), .C(new_n579_), .Y(new_n582_));
  INVX1    g0101(.A(new_n580_), .Y(new_n583_));
  INVX1    g0102(.A(new_n535_), .Y(new_n584_));
  NOR3X1   g0103(.A(new_n562_), .B(new_n584_), .C(new_n524_), .Y(new_n585_));
  OAI22X1  g0104(.A0(new_n585_), .A1(\V174(0) ), .B0(new_n583_), .B1(new_n579_), .Y(new_n586_));
  NOR2X1   g0105(.A(new_n586_), .B(new_n582_), .Y(new_n587_));
  NOR3X1   g0106(.A(new_n580_), .B(new_n579_), .C(\V59(0) ), .Y(new_n588_));
  NOR3X1   g0107(.A(new_n562_), .B(new_n524_), .C(new_n486_), .Y(new_n589_));
  NAND2X1  g0108(.A(new_n584_), .B(\V234(0) ), .Y(new_n590_));
  NAND2X1  g0109(.A(new_n535_), .B(\V194(0) ), .Y(new_n591_));
  MX2X1    g0110(.A(new_n591_), .B(new_n590_), .S0(new_n589_), .Y(new_n592_));
  OR4X1    g0111(.A(new_n592_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n593_));
  INVX1    g0112(.A(\V257(7) ), .Y(V657));
  INVX1    g0113(.A(new_n578_), .Y(new_n595_));
  INVX1    g0114(.A(new_n587_), .Y(new_n596_));
  OR4X1    g0115(.A(new_n588_), .B(new_n596_), .C(new_n595_), .D(V657), .Y(new_n597_));
  NOR4X1   g0116(.A(new_n580_), .B(new_n579_), .C(new_n496_), .D(\V59(0) ), .Y(new_n598_));
  NAND4X1  g0117(.A(new_n598_), .B(new_n587_), .C(new_n577_), .D(new_n576_), .Y(new_n599_));
  NAND3X1  g0118(.A(new_n599_), .B(new_n597_), .C(new_n593_), .Y(new_n600_));
  NOR3X1   g0119(.A(\V60(0) ), .B(\V59(0) ), .C(\V56(0) ), .Y(new_n601_));
  NOR3X1   g0120(.A(new_n601_), .B(new_n510_), .C(\V292(0) ), .Y(new_n602_));
  MX2X1    g0121(.A(\V32(5) ), .B(\V32(2) ), .S0(new_n602_), .Y(new_n603_));
  MX2X1    g0122(.A(new_n603_), .B(new_n600_), .S0(new_n575_), .Y(new_n604_));
  INVX1    g0123(.A(\V60(0) ), .Y(new_n605_));
  INVX1    g0124(.A(new_n562_), .Y(new_n606_));
  AOI21X1  g0125(.A0(new_n606_), .A1(new_n559_), .B0(new_n605_), .Y(new_n607_));
  AOI21X1  g0126(.A0(new_n570_), .A1(new_n526_), .B0(new_n607_), .Y(new_n608_));
  INVX1    g0127(.A(new_n608_), .Y(new_n609_));
  AND2X1   g0128(.A(new_n609_), .B(new_n604_), .Y(new_n610_));
  AND2X1   g0129(.A(new_n608_), .B(\V78(4) ), .Y(new_n611_));
  MX2X1    g0130(.A(new_n611_), .B(new_n610_), .S0(new_n571_), .Y(\V1243(0) ));
  INVX1    g0131(.A(\V1243(0) ), .Y(\V321(2) ));
  AND2X1   g0132(.A(\V288(1) ), .B(\V288(0) ), .Y(new_n614_));
  INVX1    g0133(.A(\V288(0) ), .Y(new_n615_));
  AND2X1   g0134(.A(\V288(1) ), .B(new_n615_), .Y(new_n616_));
  INVX1    g0135(.A(new_n616_), .Y(new_n617_));
  INVX1    g0136(.A(\V288(2) ), .Y(new_n618_));
  AND2X1   g0137(.A(\V288(3) ), .B(new_n618_), .Y(new_n619_));
  INVX1    g0138(.A(\V288(4) ), .Y(new_n620_));
  AND2X1   g0139(.A(\V288(5) ), .B(new_n620_), .Y(new_n621_));
  INVX1    g0140(.A(\V288(6) ), .Y(new_n622_));
  AND2X1   g0141(.A(\V288(7) ), .B(new_n622_), .Y(new_n623_));
  XOR2X1   g0142(.A(new_n623_), .B(new_n621_), .Y(new_n624_));
  XOR2X1   g0143(.A(new_n624_), .B(new_n619_), .Y(new_n625_));
  XOR2X1   g0144(.A(new_n625_), .B(new_n617_), .Y(new_n626_));
  OR2X1    g0145(.A(new_n625_), .B(new_n617_), .Y(new_n627_));
  INVX1    g0146(.A(\V288(1) ), .Y(new_n628_));
  AND2X1   g0147(.A(new_n628_), .B(\V288(0) ), .Y(new_n629_));
  INVX1    g0148(.A(\V288(3) ), .Y(new_n630_));
  AND2X1   g0149(.A(new_n630_), .B(\V288(2) ), .Y(new_n631_));
  OR2X1    g0150(.A(\V288(5) ), .B(new_n620_), .Y(new_n632_));
  XOR2X1   g0151(.A(\V288(7) ), .B(new_n622_), .Y(new_n633_));
  XOR2X1   g0152(.A(new_n633_), .B(new_n632_), .Y(new_n634_));
  INVX1    g0153(.A(\V288(5) ), .Y(new_n635_));
  OR2X1    g0154(.A(new_n635_), .B(\V288(4) ), .Y(new_n636_));
  NOR2X1   g0155(.A(new_n623_), .B(new_n636_), .Y(new_n637_));
  XOR2X1   g0156(.A(new_n637_), .B(new_n634_), .Y(new_n638_));
  XOR2X1   g0157(.A(new_n638_), .B(new_n631_), .Y(new_n639_));
  XOR2X1   g0158(.A(new_n623_), .B(new_n636_), .Y(new_n640_));
  AND2X1   g0159(.A(new_n640_), .B(new_n619_), .Y(new_n641_));
  XOR2X1   g0160(.A(new_n641_), .B(new_n639_), .Y(new_n642_));
  XOR2X1   g0161(.A(new_n642_), .B(new_n629_), .Y(new_n643_));
  XOR2X1   g0162(.A(new_n643_), .B(new_n627_), .Y(new_n644_));
  XOR2X1   g0163(.A(new_n644_), .B(new_n626_), .Y(new_n645_));
  NAND2X1  g0164(.A(new_n584_), .B(\V223(2) ), .Y(new_n646_));
  NAND2X1  g0165(.A(new_n535_), .B(\V183(2) ), .Y(new_n647_));
  MX2X1    g0166(.A(new_n647_), .B(new_n646_), .S0(new_n589_), .Y(new_n648_));
  OR4X1    g0167(.A(new_n648_), .B(new_n587_), .C(new_n574_), .D(new_n578_), .Y(new_n649_));
  NOR4X1   g0168(.A(new_n649_), .B(new_n608_), .C(new_n588_), .D(new_n574_), .Y(new_n650_));
  AND2X1   g0169(.A(new_n608_), .B(\V32(2) ), .Y(new_n651_));
  MX2X1    g0170(.A(new_n651_), .B(new_n650_), .S0(new_n571_), .Y(\V1213(2) ));
  XOR2X1   g0171(.A(\V1213(2) ), .B(new_n645_), .Y(new_n653_));
  NOR2X1   g0172(.A(new_n644_), .B(new_n626_), .Y(new_n654_));
  OR2X1    g0173(.A(new_n630_), .B(\V288(2) ), .Y(new_n655_));
  XOR2X1   g0174(.A(new_n624_), .B(new_n655_), .Y(new_n656_));
  AND2X1   g0175(.A(new_n656_), .B(new_n616_), .Y(new_n657_));
  OR2X1    g0176(.A(new_n624_), .B(new_n655_), .Y(new_n658_));
  XOR2X1   g0177(.A(new_n658_), .B(new_n639_), .Y(new_n659_));
  AND2X1   g0178(.A(new_n659_), .B(new_n657_), .Y(new_n660_));
  INVX1    g0179(.A(new_n629_), .Y(new_n661_));
  AOI21X1  g0180(.A0(new_n642_), .A1(new_n627_), .B0(new_n661_), .Y(new_n662_));
  OR2X1    g0181(.A(new_n662_), .B(new_n660_), .Y(new_n663_));
  OR2X1    g0182(.A(new_n623_), .B(new_n636_), .Y(new_n664_));
  XOR2X1   g0183(.A(new_n664_), .B(new_n634_), .Y(new_n665_));
  AND2X1   g0184(.A(new_n641_), .B(new_n665_), .Y(new_n666_));
  INVX1    g0185(.A(new_n631_), .Y(new_n667_));
  AOI21X1  g0186(.A0(new_n658_), .A1(new_n638_), .B0(new_n667_), .Y(new_n668_));
  OR2X1    g0187(.A(new_n668_), .B(new_n666_), .Y(new_n669_));
  AND2X1   g0188(.A(\V288(3) ), .B(\V288(2) ), .Y(new_n670_));
  INVX1    g0189(.A(\V288(7) ), .Y(new_n671_));
  AND2X1   g0190(.A(new_n671_), .B(\V288(6) ), .Y(new_n672_));
  NOR3X1   g0191(.A(new_n672_), .B(new_n623_), .C(new_n636_), .Y(new_n673_));
  NOR4X1   g0192(.A(new_n672_), .B(new_n623_), .C(\V288(5) ), .D(new_n620_), .Y(new_n674_));
  OR2X1    g0193(.A(new_n674_), .B(new_n673_), .Y(new_n675_));
  NAND2X1  g0194(.A(\V288(5) ), .B(\V288(4) ), .Y(new_n676_));
  NOR2X1   g0195(.A(\V288(7) ), .B(\V288(6) ), .Y(new_n677_));
  XOR2X1   g0196(.A(new_n677_), .B(new_n676_), .Y(new_n678_));
  XOR2X1   g0197(.A(new_n678_), .B(new_n675_), .Y(new_n679_));
  XOR2X1   g0198(.A(new_n679_), .B(new_n670_), .Y(new_n680_));
  XOR2X1   g0199(.A(new_n680_), .B(new_n669_), .Y(new_n681_));
  XOR2X1   g0200(.A(new_n681_), .B(new_n614_), .Y(new_n682_));
  XOR2X1   g0201(.A(new_n682_), .B(new_n663_), .Y(new_n683_));
  AND2X1   g0202(.A(new_n683_), .B(new_n654_), .Y(new_n684_));
  OR4X1    g0203(.A(\V288(5) ), .B(\V288(4) ), .C(\V288(7) ), .D(\V288(6) ), .Y(new_n685_));
  INVX1    g0204(.A(new_n679_), .Y(new_n686_));
  NOR2X1   g0205(.A(new_n668_), .B(new_n666_), .Y(new_n687_));
  INVX1    g0206(.A(new_n670_), .Y(new_n688_));
  AOI21X1  g0207(.A0(new_n679_), .A1(new_n687_), .B0(new_n688_), .Y(new_n689_));
  AOI21X1  g0208(.A0(new_n686_), .A1(new_n669_), .B0(new_n689_), .Y(new_n690_));
  XOR2X1   g0209(.A(new_n690_), .B(new_n685_), .Y(new_n691_));
  XOR2X1   g0210(.A(new_n680_), .B(new_n687_), .Y(new_n692_));
  INVX1    g0211(.A(new_n614_), .Y(new_n693_));
  OR4X1    g0212(.A(new_n642_), .B(new_n627_), .C(new_n628_), .D(new_n615_), .Y(new_n694_));
  OAI21X1  g0213(.A0(new_n681_), .A1(new_n693_), .B0(new_n694_), .Y(new_n695_));
  AOI21X1  g0214(.A0(new_n692_), .A1(new_n663_), .B0(new_n695_), .Y(new_n696_));
  XOR2X1   g0215(.A(new_n696_), .B(new_n691_), .Y(new_n697_));
  XOR2X1   g0216(.A(new_n697_), .B(new_n684_), .Y(new_n698_));
  NAND2X1  g0217(.A(new_n584_), .B(\V223(0) ), .Y(new_n699_));
  NAND2X1  g0218(.A(new_n535_), .B(\V183(0) ), .Y(new_n700_));
  MX2X1    g0219(.A(new_n700_), .B(new_n699_), .S0(new_n589_), .Y(new_n701_));
  OR4X1    g0220(.A(new_n701_), .B(new_n587_), .C(new_n574_), .D(new_n578_), .Y(new_n702_));
  NOR4X1   g0221(.A(new_n702_), .B(new_n608_), .C(new_n588_), .D(new_n574_), .Y(new_n703_));
  INVX1    g0222(.A(\V32(0) ), .Y(new_n704_));
  NOR3X1   g0223(.A(new_n607_), .B(new_n571_), .C(new_n704_), .Y(new_n705_));
  AOI21X1  g0224(.A0(new_n703_), .A1(new_n571_), .B0(new_n705_), .Y(new_n706_));
  XOR2X1   g0225(.A(new_n706_), .B(new_n698_), .Y(new_n707_));
  XOR2X1   g0226(.A(new_n683_), .B(new_n654_), .Y(new_n708_));
  NAND2X1  g0227(.A(new_n584_), .B(\V223(1) ), .Y(new_n709_));
  NAND2X1  g0228(.A(new_n535_), .B(\V183(1) ), .Y(new_n710_));
  MX2X1    g0229(.A(new_n710_), .B(new_n709_), .S0(new_n589_), .Y(new_n711_));
  OR4X1    g0230(.A(new_n711_), .B(new_n587_), .C(new_n574_), .D(new_n578_), .Y(new_n712_));
  NOR4X1   g0231(.A(new_n712_), .B(new_n608_), .C(new_n588_), .D(new_n574_), .Y(new_n713_));
  INVX1    g0232(.A(\V32(1) ), .Y(new_n714_));
  NOR3X1   g0233(.A(new_n607_), .B(new_n571_), .C(new_n714_), .Y(new_n715_));
  AOI21X1  g0234(.A0(new_n713_), .A1(new_n571_), .B0(new_n715_), .Y(new_n716_));
  XOR2X1   g0235(.A(new_n716_), .B(new_n708_), .Y(new_n717_));
  NAND3X1  g0236(.A(\V149(3) ), .B(new_n527_), .C(new_n501_), .Y(new_n718_));
  NOR4X1   g0237(.A(new_n718_), .B(new_n498_), .C(\V149(4) ), .D(\V149(6) ), .Y(new_n719_));
  AND2X1   g0238(.A(new_n719_), .B(new_n493_), .Y(new_n720_));
  NAND2X1  g0239(.A(new_n584_), .B(\V223(3) ), .Y(new_n721_));
  NAND2X1  g0240(.A(new_n535_), .B(\V183(3) ), .Y(new_n722_));
  MX2X1    g0241(.A(new_n722_), .B(new_n721_), .S0(new_n589_), .Y(new_n723_));
  OR4X1    g0242(.A(new_n723_), .B(new_n587_), .C(new_n574_), .D(new_n578_), .Y(new_n724_));
  NOR4X1   g0243(.A(new_n724_), .B(new_n608_), .C(new_n588_), .D(new_n574_), .Y(new_n725_));
  INVX1    g0244(.A(\V32(3) ), .Y(new_n726_));
  NOR3X1   g0245(.A(new_n607_), .B(new_n571_), .C(new_n726_), .Y(new_n727_));
  AOI21X1  g0246(.A0(new_n725_), .A1(new_n571_), .B0(new_n727_), .Y(new_n728_));
  XOR2X1   g0247(.A(new_n728_), .B(new_n626_), .Y(new_n729_));
  NOR4X1   g0248(.A(new_n729_), .B(new_n720_), .C(new_n717_), .D(new_n707_), .Y(new_n730_));
  NAND3X1  g0249(.A(new_n730_), .B(new_n653_), .C(new_n614_), .Y(new_n731_));
  INVX1    g0250(.A(new_n731_), .Y(new_n732_));
  INVX1    g0251(.A(\V32(2) ), .Y(new_n733_));
  NOR3X1   g0252(.A(new_n607_), .B(new_n571_), .C(new_n733_), .Y(new_n734_));
  AOI21X1  g0253(.A0(new_n650_), .A1(new_n571_), .B0(new_n734_), .Y(new_n735_));
  XOR2X1   g0254(.A(new_n642_), .B(new_n625_), .Y(new_n736_));
  XOR2X1   g0255(.A(new_n736_), .B(new_n735_), .Y(new_n737_));
  INVX1    g0256(.A(new_n685_), .Y(new_n738_));
  XOR2X1   g0257(.A(new_n690_), .B(new_n738_), .Y(new_n739_));
  AND2X1   g0258(.A(new_n642_), .B(new_n625_), .Y(new_n740_));
  AND2X1   g0259(.A(new_n740_), .B(new_n681_), .Y(new_n741_));
  XOR2X1   g0260(.A(new_n741_), .B(new_n739_), .Y(new_n742_));
  XOR2X1   g0261(.A(new_n742_), .B(new_n706_), .Y(new_n743_));
  XOR2X1   g0262(.A(new_n740_), .B(new_n681_), .Y(new_n744_));
  XOR2X1   g0263(.A(new_n744_), .B(new_n716_), .Y(new_n745_));
  XOR2X1   g0264(.A(new_n728_), .B(new_n656_), .Y(new_n746_));
  OR4X1    g0265(.A(new_n746_), .B(new_n745_), .C(new_n743_), .D(new_n720_), .Y(new_n747_));
  NOR3X1   g0266(.A(new_n747_), .B(new_n737_), .C(new_n688_), .Y(new_n748_));
  XOR2X1   g0267(.A(new_n638_), .B(new_n624_), .Y(new_n749_));
  XOR2X1   g0268(.A(new_n749_), .B(new_n735_), .Y(new_n750_));
  AND2X1   g0269(.A(new_n638_), .B(new_n624_), .Y(new_n751_));
  AND2X1   g0270(.A(new_n751_), .B(new_n679_), .Y(new_n752_));
  XOR2X1   g0271(.A(new_n752_), .B(new_n685_), .Y(new_n753_));
  XOR2X1   g0272(.A(new_n753_), .B(new_n706_), .Y(new_n754_));
  XOR2X1   g0273(.A(new_n751_), .B(new_n679_), .Y(new_n755_));
  XOR2X1   g0274(.A(new_n755_), .B(new_n716_), .Y(new_n756_));
  XOR2X1   g0275(.A(new_n728_), .B(new_n640_), .Y(new_n757_));
  OR4X1    g0276(.A(new_n757_), .B(new_n756_), .C(new_n754_), .D(new_n720_), .Y(new_n758_));
  NOR3X1   g0277(.A(new_n758_), .B(new_n750_), .C(new_n676_), .Y(new_n759_));
  AND2X1   g0278(.A(new_n608_), .B(\V32(3) ), .Y(new_n760_));
  MX2X1    g0279(.A(new_n760_), .B(new_n725_), .S0(new_n571_), .Y(\V1213(3) ));
  AND2X1   g0280(.A(new_n608_), .B(\V32(0) ), .Y(new_n762_));
  MX2X1    g0281(.A(new_n762_), .B(new_n703_), .S0(new_n571_), .Y(\V1213(0) ));
  AND2X1   g0282(.A(new_n608_), .B(\V32(1) ), .Y(new_n764_));
  MX2X1    g0283(.A(new_n764_), .B(new_n713_), .S0(new_n571_), .Y(\V1213(1) ));
  OR4X1    g0284(.A(new_n720_), .B(\V1213(1) ), .C(\V1213(0) ), .D(new_n735_), .Y(new_n766_));
  NOR4X1   g0285(.A(new_n766_), .B(\V1213(3) ), .C(new_n671_), .D(new_n622_), .Y(new_n767_));
  INVX1    g0286(.A(new_n677_), .Y(new_n768_));
  NOR4X1   g0287(.A(\V1213(3) ), .B(new_n720_), .C(\V1213(1) ), .D(\V1213(0) ), .Y(new_n769_));
  NAND3X1  g0288(.A(new_n769_), .B(new_n768_), .C(new_n735_), .Y(new_n770_));
  INVX1    g0289(.A(new_n770_), .Y(new_n771_));
  NOR2X1   g0290(.A(\V288(5) ), .B(\V288(4) ), .Y(new_n772_));
  OR2X1    g0291(.A(\V288(7) ), .B(new_n622_), .Y(new_n773_));
  XOR2X1   g0292(.A(new_n773_), .B(new_n735_), .Y(new_n774_));
  OAI21X1  g0293(.A0(new_n671_), .A1(new_n622_), .B0(new_n620_), .Y(new_n775_));
  MX2X1    g0294(.A(new_n775_), .B(new_n685_), .S0(new_n621_), .Y(new_n776_));
  XOR2X1   g0295(.A(new_n776_), .B(new_n706_), .Y(new_n777_));
  NOR4X1   g0296(.A(new_n635_), .B(\V288(4) ), .C(\V288(7) ), .D(new_n622_), .Y(new_n778_));
  INVX1    g0297(.A(new_n632_), .Y(new_n779_));
  AND2X1   g0298(.A(new_n638_), .B(new_n640_), .Y(new_n780_));
  XOR2X1   g0299(.A(new_n780_), .B(new_n755_), .Y(new_n781_));
  MX2X1    g0300(.A(new_n781_), .B(new_n679_), .S0(new_n779_), .Y(new_n782_));
  XOR2X1   g0301(.A(new_n782_), .B(new_n778_), .Y(new_n783_));
  MX2X1    g0302(.A(new_n783_), .B(new_n679_), .S0(new_n621_), .Y(new_n784_));
  XOR2X1   g0303(.A(new_n784_), .B(new_n716_), .Y(new_n785_));
  OR2X1    g0304(.A(new_n671_), .B(\V288(6) ), .Y(new_n786_));
  XOR2X1   g0305(.A(new_n786_), .B(new_n728_), .Y(new_n787_));
  OR4X1    g0306(.A(new_n787_), .B(new_n785_), .C(new_n777_), .D(new_n720_), .Y(new_n788_));
  NOR3X1   g0307(.A(new_n788_), .B(new_n774_), .C(new_n772_), .Y(new_n789_));
  NOR2X1   g0308(.A(\V288(3) ), .B(\V288(2) ), .Y(new_n790_));
  XOR2X1   g0309(.A(new_n624_), .B(new_n619_), .Y(new_n791_));
  XOR2X1   g0310(.A(new_n736_), .B(new_n656_), .Y(new_n792_));
  MX2X1    g0311(.A(new_n792_), .B(new_n642_), .S0(new_n631_), .Y(new_n793_));
  XOR2X1   g0312(.A(new_n793_), .B(new_n791_), .Y(new_n794_));
  MX2X1    g0313(.A(new_n794_), .B(new_n642_), .S0(new_n619_), .Y(new_n795_));
  XOR2X1   g0314(.A(new_n795_), .B(new_n735_), .Y(new_n796_));
  AND2X1   g0315(.A(new_n793_), .B(new_n791_), .Y(new_n797_));
  AND2X1   g0316(.A(new_n642_), .B(new_n656_), .Y(new_n798_));
  XOR2X1   g0317(.A(new_n798_), .B(new_n744_), .Y(new_n799_));
  MX2X1    g0318(.A(new_n799_), .B(new_n681_), .S0(new_n631_), .Y(new_n800_));
  AND2X1   g0319(.A(new_n800_), .B(new_n797_), .Y(new_n801_));
  NOR3X1   g0320(.A(new_n692_), .B(new_n659_), .C(new_n625_), .Y(new_n802_));
  XOR2X1   g0321(.A(new_n802_), .B(new_n742_), .Y(new_n803_));
  MX2X1    g0322(.A(new_n803_), .B(new_n739_), .S0(new_n631_), .Y(new_n804_));
  XOR2X1   g0323(.A(new_n804_), .B(new_n801_), .Y(new_n805_));
  MX2X1    g0324(.A(new_n805_), .B(new_n739_), .S0(new_n619_), .Y(new_n806_));
  XOR2X1   g0325(.A(new_n806_), .B(new_n706_), .Y(new_n807_));
  INVX1    g0326(.A(new_n720_), .Y(new_n808_));
  XOR2X1   g0327(.A(new_n800_), .B(new_n797_), .Y(new_n809_));
  MX2X1    g0328(.A(new_n809_), .B(new_n681_), .S0(new_n619_), .Y(new_n810_));
  XOR2X1   g0329(.A(new_n810_), .B(\V1213(1) ), .Y(new_n811_));
  XOR2X1   g0330(.A(new_n625_), .B(new_n655_), .Y(new_n812_));
  XOR2X1   g0331(.A(new_n812_), .B(\V1213(3) ), .Y(new_n813_));
  NAND3X1  g0332(.A(new_n813_), .B(new_n811_), .C(new_n808_), .Y(new_n814_));
  OR4X1    g0333(.A(new_n814_), .B(new_n807_), .C(new_n796_), .D(new_n790_), .Y(new_n815_));
  INVX1    g0334(.A(new_n815_), .Y(new_n816_));
  NOR2X1   g0335(.A(\V288(1) ), .B(\V288(0) ), .Y(new_n817_));
  XOR2X1   g0336(.A(new_n643_), .B(new_n657_), .Y(new_n818_));
  XOR2X1   g0337(.A(new_n625_), .B(new_n616_), .Y(new_n819_));
  XOR2X1   g0338(.A(new_n645_), .B(new_n626_), .Y(new_n820_));
  MX2X1    g0339(.A(new_n820_), .B(new_n818_), .S0(new_n629_), .Y(new_n821_));
  XOR2X1   g0340(.A(new_n821_), .B(new_n819_), .Y(new_n822_));
  MX2X1    g0341(.A(new_n822_), .B(new_n818_), .S0(new_n616_), .Y(new_n823_));
  XOR2X1   g0342(.A(new_n823_), .B(new_n735_), .Y(new_n824_));
  AND2X1   g0343(.A(new_n821_), .B(new_n819_), .Y(new_n825_));
  AND2X1   g0344(.A(new_n818_), .B(new_n626_), .Y(new_n826_));
  XOR2X1   g0345(.A(new_n826_), .B(new_n708_), .Y(new_n827_));
  MX2X1    g0346(.A(new_n827_), .B(new_n683_), .S0(new_n629_), .Y(new_n828_));
  AND2X1   g0347(.A(new_n828_), .B(new_n825_), .Y(new_n829_));
  INVX1    g0348(.A(new_n626_), .Y(new_n830_));
  NOR2X1   g0349(.A(new_n662_), .B(new_n660_), .Y(new_n831_));
  XOR2X1   g0350(.A(new_n682_), .B(new_n831_), .Y(new_n832_));
  NOR3X1   g0351(.A(new_n832_), .B(new_n644_), .C(new_n830_), .Y(new_n833_));
  XOR2X1   g0352(.A(new_n833_), .B(new_n698_), .Y(new_n834_));
  MX2X1    g0353(.A(new_n834_), .B(new_n697_), .S0(new_n629_), .Y(new_n835_));
  XOR2X1   g0354(.A(new_n835_), .B(new_n829_), .Y(new_n836_));
  MX2X1    g0355(.A(new_n836_), .B(new_n697_), .S0(new_n616_), .Y(new_n837_));
  XOR2X1   g0356(.A(new_n837_), .B(new_n706_), .Y(new_n838_));
  XOR2X1   g0357(.A(new_n828_), .B(new_n825_), .Y(new_n839_));
  MX2X1    g0358(.A(new_n839_), .B(new_n683_), .S0(new_n616_), .Y(new_n840_));
  XOR2X1   g0359(.A(new_n840_), .B(\V1213(1) ), .Y(new_n841_));
  XOR2X1   g0360(.A(new_n626_), .B(new_n616_), .Y(new_n842_));
  XOR2X1   g0361(.A(new_n842_), .B(\V1213(3) ), .Y(new_n843_));
  NAND3X1  g0362(.A(new_n843_), .B(new_n841_), .C(new_n808_), .Y(new_n844_));
  NOR4X1   g0363(.A(new_n844_), .B(new_n838_), .C(new_n824_), .D(new_n817_), .Y(new_n845_));
  OR4X1    g0364(.A(new_n845_), .B(new_n816_), .C(new_n720_), .D(new_n578_), .Y(new_n846_));
  OR4X1    g0365(.A(new_n846_), .B(new_n789_), .C(new_n771_), .D(new_n767_), .Y(new_n847_));
  NOR4X1   g0366(.A(new_n847_), .B(new_n759_), .C(new_n748_), .D(new_n732_), .Y(V356));
  XOR2X1   g0367(.A(new_n735_), .B(new_n818_), .Y(new_n849_));
  XOR2X1   g0368(.A(new_n706_), .B(new_n697_), .Y(new_n850_));
  XOR2X1   g0369(.A(new_n716_), .B(new_n683_), .Y(new_n851_));
  XOR2X1   g0370(.A(new_n728_), .B(new_n830_), .Y(new_n852_));
  OR4X1    g0371(.A(new_n852_), .B(new_n851_), .C(new_n850_), .D(new_n720_), .Y(new_n853_));
  NOR3X1   g0372(.A(new_n853_), .B(new_n849_), .C(new_n693_), .Y(new_n854_));
  XOR2X1   g0373(.A(new_n735_), .B(new_n642_), .Y(new_n855_));
  XOR2X1   g0374(.A(new_n706_), .B(new_n739_), .Y(new_n856_));
  XOR2X1   g0375(.A(new_n716_), .B(new_n681_), .Y(new_n857_));
  XOR2X1   g0376(.A(new_n728_), .B(new_n625_), .Y(new_n858_));
  OR4X1    g0377(.A(new_n858_), .B(new_n857_), .C(new_n856_), .D(new_n720_), .Y(new_n859_));
  NOR3X1   g0378(.A(new_n859_), .B(new_n855_), .C(new_n688_), .Y(new_n860_));
  XOR2X1   g0379(.A(new_n735_), .B(new_n638_), .Y(new_n861_));
  XOR2X1   g0380(.A(new_n706_), .B(new_n685_), .Y(new_n862_));
  XOR2X1   g0381(.A(new_n716_), .B(new_n679_), .Y(new_n863_));
  XOR2X1   g0382(.A(new_n728_), .B(new_n624_), .Y(new_n864_));
  OR4X1    g0383(.A(new_n864_), .B(new_n863_), .C(new_n862_), .D(new_n720_), .Y(new_n865_));
  NOR3X1   g0384(.A(new_n865_), .B(new_n861_), .C(new_n676_), .Y(new_n866_));
  OR4X1    g0385(.A(new_n720_), .B(\V1213(1) ), .C(\V1213(0) ), .D(new_n735_), .Y(new_n867_));
  NOR4X1   g0386(.A(new_n867_), .B(new_n728_), .C(new_n671_), .D(new_n622_), .Y(new_n868_));
  NOR4X1   g0387(.A(new_n728_), .B(new_n720_), .C(\V1213(1) ), .D(\V1213(0) ), .Y(new_n869_));
  NAND3X1  g0388(.A(new_n869_), .B(new_n735_), .C(\V288(6) ), .Y(new_n870_));
  INVX1    g0389(.A(new_n870_), .Y(new_n871_));
  XOR2X1   g0390(.A(new_n749_), .B(new_n640_), .Y(new_n872_));
  MX2X1    g0391(.A(new_n872_), .B(new_n638_), .S0(new_n779_), .Y(new_n873_));
  XOR2X1   g0392(.A(new_n873_), .B(new_n735_), .Y(new_n874_));
  AND2X1   g0393(.A(new_n780_), .B(new_n755_), .Y(new_n875_));
  XOR2X1   g0394(.A(new_n875_), .B(new_n753_), .Y(new_n876_));
  MX2X1    g0395(.A(new_n876_), .B(new_n685_), .S0(new_n779_), .Y(new_n877_));
  XOR2X1   g0396(.A(new_n877_), .B(new_n706_), .Y(new_n878_));
  XOR2X1   g0397(.A(new_n782_), .B(new_n716_), .Y(new_n879_));
  XOR2X1   g0398(.A(new_n623_), .B(new_n621_), .Y(new_n880_));
  XOR2X1   g0399(.A(new_n880_), .B(new_n728_), .Y(new_n881_));
  OR4X1    g0400(.A(new_n881_), .B(new_n879_), .C(new_n878_), .D(new_n720_), .Y(new_n882_));
  NOR3X1   g0401(.A(new_n882_), .B(new_n874_), .C(new_n620_), .Y(new_n883_));
  XOR2X1   g0402(.A(new_n793_), .B(\V1213(2) ), .Y(new_n884_));
  XOR2X1   g0403(.A(new_n804_), .B(new_n706_), .Y(new_n885_));
  XOR2X1   g0404(.A(new_n800_), .B(new_n716_), .Y(new_n886_));
  XOR2X1   g0405(.A(new_n791_), .B(new_n728_), .Y(new_n887_));
  NOR4X1   g0406(.A(new_n887_), .B(new_n886_), .C(new_n885_), .D(new_n720_), .Y(new_n888_));
  NAND3X1  g0407(.A(new_n888_), .B(new_n884_), .C(\V288(2) ), .Y(new_n889_));
  INVX1    g0408(.A(new_n889_), .Y(new_n890_));
  XOR2X1   g0409(.A(new_n821_), .B(new_n735_), .Y(new_n891_));
  XOR2X1   g0410(.A(new_n835_), .B(new_n706_), .Y(new_n892_));
  XOR2X1   g0411(.A(new_n828_), .B(\V1213(1) ), .Y(new_n893_));
  XOR2X1   g0412(.A(new_n819_), .B(\V1213(3) ), .Y(new_n894_));
  NAND3X1  g0413(.A(new_n894_), .B(new_n893_), .C(new_n808_), .Y(new_n895_));
  NOR4X1   g0414(.A(new_n895_), .B(new_n892_), .C(new_n891_), .D(new_n615_), .Y(new_n896_));
  OR4X1    g0415(.A(new_n896_), .B(new_n890_), .C(new_n883_), .D(new_n578_), .Y(new_n897_));
  OR4X1    g0416(.A(new_n897_), .B(new_n871_), .C(new_n868_), .D(new_n866_), .Y(new_n898_));
  NOR3X1   g0417(.A(new_n898_), .B(new_n860_), .C(new_n854_), .Y(V357));
  AND2X1   g0418(.A(\V13(0) ), .B(\V10(0) ), .Y(V373));
  AND2X1   g0419(.A(\V9(0) ), .B(\V1(0) ), .Y(V1423));
  AND2X1   g0420(.A(\V2(0) ), .B(\V9(0) ), .Y(V1258));
  AND2X1   g0421(.A(\V9(0) ), .B(\V7(0) ), .Y(V787));
  INVX1    g0422(.A(\V13(0) ), .Y(new_n904_));
  AND2X1   g0423(.A(\V109(0) ), .B(new_n904_), .Y(new_n905_));
  NOR3X1   g0424(.A(V787), .B(V1258), .C(V1423), .Y(new_n906_));
  AND2X1   g0425(.A(\V5(0) ), .B(\V9(0) ), .Y(V778));
  AND2X1   g0426(.A(\V8(0) ), .B(\V9(0) ), .Y(V1387));
  AND2X1   g0427(.A(\V6(0) ), .B(\V9(0) ), .Y(V780));
  NOR3X1   g0428(.A(V780), .B(V1387), .C(V778), .Y(new_n910_));
  AND2X1   g0429(.A(\V71(0) ), .B(\V202(0) ), .Y(new_n911_));
  AND2X1   g0430(.A(new_n911_), .B(new_n904_), .Y(new_n912_));
  OAI21X1  g0431(.A0(\V3(0) ), .A1(\V4(0) ), .B0(\V9(0) ), .Y(new_n913_));
  NAND3X1  g0432(.A(new_n913_), .B(new_n910_), .C(new_n906_), .Y(\V375(0) ));
  NAND2X1  g0433(.A(\V165(1) ), .B(\V203(0) ), .Y(new_n915_));
  NOR3X1   g0434(.A(new_n915_), .B(new_n512_), .C(\V165(0) ), .Y(new_n916_));
  OR2X1    g0435(.A(new_n916_), .B(\V35(0) ), .Y(new_n917_));
  AND2X1   g0436(.A(new_n917_), .B(\V203(0) ), .Y(V377));
  INVX1    g0437(.A(\V240(0) ), .Y(new_n919_));
  NOR3X1   g0438(.A(new_n513_), .B(\V165(2) ), .C(new_n511_), .Y(new_n920_));
  NOR3X1   g0439(.A(new_n920_), .B(new_n919_), .C(\V172(0) ), .Y(V1719));
  INVX1    g0440(.A(V1719), .Y(new_n922_));
  INVX1    g0441(.A(\V194(4) ), .Y(new_n923_));
  INVX1    g0442(.A(\V194(2) ), .Y(new_n924_));
  INVX1    g0443(.A(\V194(1) ), .Y(new_n925_));
  NAND4X1  g0444(.A(\V194(3) ), .B(\V199(0) ), .C(\V199(2) ), .D(\V199(4) ), .Y(new_n926_));
  NOR4X1   g0445(.A(new_n926_), .B(new_n925_), .C(new_n924_), .D(new_n923_), .Y(new_n927_));
  NAND3X1  g0446(.A(new_n927_), .B(\V199(1) ), .C(\V199(3) ), .Y(new_n928_));
  NOR3X1   g0447(.A(new_n928_), .B(new_n922_), .C(\V248(0) ), .Y(new_n929_));
  INVX1    g0448(.A(\V247(0) ), .Y(new_n930_));
  NAND4X1  g0449(.A(\V246(0) ), .B(\V245(0) ), .C(\V244(0) ), .D(\V243(0) ), .Y(new_n931_));
  NOR4X1   g0450(.A(new_n931_), .B(new_n922_), .C(new_n930_), .D(\V248(0) ), .Y(new_n932_));
  INVX1    g0451(.A(\V239(4) ), .Y(new_n933_));
  OR2X1    g0452(.A(new_n535_), .B(new_n933_), .Y(new_n934_));
  NAND2X1  g0453(.A(new_n535_), .B(\V199(4) ), .Y(new_n935_));
  MX2X1    g0454(.A(new_n935_), .B(new_n934_), .S0(new_n589_), .Y(new_n936_));
  NOR4X1   g0455(.A(new_n936_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n937_));
  INVX1    g0456(.A(\V32(11) ), .Y(new_n938_));
  INVX1    g0457(.A(new_n602_), .Y(new_n939_));
  NOR3X1   g0458(.A(new_n939_), .B(new_n575_), .C(new_n938_), .Y(new_n940_));
  MX2X1    g0459(.A(new_n940_), .B(new_n937_), .S0(new_n575_), .Y(new_n941_));
  AND2X1   g0460(.A(new_n941_), .B(new_n609_), .Y(new_n942_));
  AND2X1   g0461(.A(new_n608_), .B(\V88(1) ), .Y(new_n943_));
  MX2X1    g0462(.A(new_n943_), .B(new_n942_), .S0(new_n571_), .Y(\V1243(9) ));
  INVX1    g0463(.A(\V1243(9) ), .Y(new_n945_));
  NAND2X1  g0464(.A(new_n584_), .B(\V239(2) ), .Y(new_n946_));
  NAND2X1  g0465(.A(new_n535_), .B(\V199(2) ), .Y(new_n947_));
  MX2X1    g0466(.A(new_n947_), .B(new_n946_), .S0(new_n589_), .Y(new_n948_));
  NOR4X1   g0467(.A(new_n948_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n949_));
  INVX1    g0468(.A(\V32(9) ), .Y(new_n950_));
  NOR3X1   g0469(.A(new_n939_), .B(new_n575_), .C(new_n950_), .Y(new_n951_));
  MX2X1    g0470(.A(new_n951_), .B(new_n949_), .S0(new_n575_), .Y(new_n952_));
  AND2X1   g0471(.A(new_n952_), .B(new_n609_), .Y(new_n953_));
  AND2X1   g0472(.A(new_n608_), .B(\V84(5) ), .Y(new_n954_));
  MX2X1    g0473(.A(new_n954_), .B(new_n953_), .S0(new_n571_), .Y(\V1243(7) ));
  INVX1    g0474(.A(\V1243(7) ), .Y(new_n956_));
  NAND2X1  g0475(.A(new_n584_), .B(\V239(3) ), .Y(new_n957_));
  NAND2X1  g0476(.A(new_n535_), .B(\V199(3) ), .Y(new_n958_));
  MX2X1    g0477(.A(new_n958_), .B(new_n957_), .S0(new_n589_), .Y(new_n959_));
  NOR4X1   g0478(.A(new_n959_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n960_));
  INVX1    g0479(.A(\V32(10) ), .Y(new_n961_));
  NOR3X1   g0480(.A(new_n939_), .B(new_n575_), .C(new_n961_), .Y(new_n962_));
  MX2X1    g0481(.A(new_n962_), .B(new_n960_), .S0(new_n575_), .Y(new_n963_));
  AND2X1   g0482(.A(new_n963_), .B(new_n609_), .Y(new_n964_));
  AND2X1   g0483(.A(new_n608_), .B(\V88(0) ), .Y(new_n965_));
  MX2X1    g0484(.A(new_n965_), .B(new_n964_), .S0(new_n571_), .Y(\V1243(8) ));
  INVX1    g0485(.A(\V1243(8) ), .Y(new_n967_));
  NOR3X1   g0486(.A(new_n896_), .B(new_n845_), .C(new_n578_), .Y(new_n968_));
  NOR3X1   g0487(.A(new_n854_), .B(new_n732_), .C(new_n578_), .Y(new_n969_));
  AOI21X1  g0488(.A0(new_n969_), .A1(new_n968_), .B0(new_n693_), .Y(new_n970_));
  NOR3X1   g0489(.A(new_n883_), .B(new_n789_), .C(new_n578_), .Y(new_n971_));
  NOR3X1   g0490(.A(new_n866_), .B(new_n759_), .C(new_n578_), .Y(new_n972_));
  AOI21X1  g0491(.A0(new_n972_), .A1(new_n971_), .B0(new_n676_), .Y(new_n973_));
  NAND3X1  g0492(.A(new_n870_), .B(new_n770_), .C(new_n595_), .Y(new_n974_));
  OR4X1    g0493(.A(new_n974_), .B(new_n868_), .C(new_n767_), .D(new_n578_), .Y(new_n975_));
  NAND3X1  g0494(.A(new_n975_), .B(\V288(7) ), .C(\V288(6) ), .Y(new_n976_));
  NAND3X1  g0495(.A(new_n889_), .B(new_n815_), .C(new_n595_), .Y(new_n977_));
  NOR4X1   g0496(.A(new_n977_), .B(new_n860_), .C(new_n748_), .D(new_n578_), .Y(new_n978_));
  OAI21X1  g0497(.A0(new_n978_), .A1(new_n688_), .B0(new_n976_), .Y(new_n979_));
  NOR3X1   g0498(.A(new_n979_), .B(new_n973_), .C(new_n970_), .Y(new_n980_));
  OR4X1    g0499(.A(new_n980_), .B(new_n967_), .C(new_n956_), .D(\V248(0) ), .Y(new_n981_));
  NOR3X1   g0500(.A(new_n981_), .B(new_n945_), .C(new_n922_), .Y(new_n982_));
  OR2X1    g0501(.A(new_n982_), .B(new_n932_), .Y(new_n983_));
  OR2X1    g0502(.A(new_n983_), .B(new_n929_), .Y(\V393(0) ));
  AND2X1   g0503(.A(V1719), .B(new_n916_), .Y(new_n985_));
  INVX1    g0504(.A(\V302(0) ), .Y(\V1864(0) ));
  NOR4X1   g0505(.A(new_n920_), .B(new_n919_), .C(\V172(0) ), .D(\V1864(0) ), .Y(new_n987_));
  NOR4X1   g0506(.A(new_n513_), .B(\V165(7) ), .C(\V165(2) ), .D(new_n511_), .Y(new_n988_));
  AND2X1   g0507(.A(new_n988_), .B(V1719), .Y(new_n989_));
  INVX1    g0508(.A(\V215(0) ), .Y(new_n990_));
  INVX1    g0509(.A(\V66(0) ), .Y(new_n991_));
  NOR4X1   g0510(.A(new_n920_), .B(new_n510_), .C(\V292(0) ), .D(new_n991_), .Y(new_n992_));
  NOR4X1   g0511(.A(new_n564_), .B(\V149(3) ), .C(new_n496_), .D(new_n527_), .Y(new_n993_));
  MX2X1    g0512(.A(new_n552_), .B(new_n546_), .S0(\V88(3) ), .Y(new_n994_));
  NOR2X1   g0513(.A(new_n994_), .B(new_n538_), .Y(new_n995_));
  OR2X1    g0514(.A(new_n995_), .B(new_n993_), .Y(new_n996_));
  OR4X1    g0515(.A(new_n996_), .B(new_n555_), .C(new_n537_), .D(\V174(0) ), .Y(new_n997_));
  AOI22X1  g0516(.A0(new_n997_), .A1(\V56(0) ), .B0(new_n992_), .B1(new_n990_), .Y(new_n998_));
  NOR3X1   g0517(.A(new_n589_), .B(new_n580_), .C(new_n493_), .Y(new_n999_));
  NOR2X1   g0518(.A(new_n999_), .B(V1719), .Y(new_n1000_));
  INVX1    g0519(.A(\V62(0) ), .Y(new_n1001_));
  NOR3X1   g0520(.A(new_n554_), .B(new_n539_), .C(new_n1001_), .Y(new_n1002_));
  AOI21X1  g0521(.A0(new_n578_), .A1(\V70(0) ), .B0(new_n1002_), .Y(new_n1003_));
  NAND4X1  g0522(.A(new_n567_), .B(new_n560_), .C(new_n558_), .D(new_n595_), .Y(new_n1004_));
  INVX1    g0523(.A(\V59(0) ), .Y(new_n1005_));
  INVX1    g0524(.A(new_n567_), .Y(new_n1006_));
  NOR2X1   g0525(.A(new_n554_), .B(new_n538_), .Y(new_n1007_));
  NOR2X1   g0526(.A(new_n994_), .B(new_n539_), .Y(new_n1008_));
  NOR3X1   g0527(.A(new_n1008_), .B(new_n1007_), .C(new_n1006_), .Y(new_n1009_));
  AOI21X1  g0528(.A0(new_n1009_), .A1(new_n595_), .B0(new_n1005_), .Y(new_n1010_));
  AOI21X1  g0529(.A0(new_n1004_), .A1(\V802(0) ), .B0(new_n1010_), .Y(new_n1011_));
  NAND4X1  g0530(.A(new_n1011_), .B(new_n1003_), .C(new_n1000_), .D(new_n998_), .Y(\V423(0) ));
  AOI21X1  g0531(.A0(V1719), .A1(\V248(0) ), .B0(\V423(0) ), .Y(new_n1013_));
  AOI21X1  g0532(.A0(new_n539_), .A1(new_n572_), .B0(new_n493_), .Y(new_n1014_));
  OR4X1    g0533(.A(new_n1014_), .B(new_n1013_), .C(\V214(0) ), .D(\V43(0) ), .Y(new_n1015_));
  OR4X1    g0534(.A(new_n1015_), .B(new_n989_), .C(new_n987_), .D(new_n929_), .Y(new_n1016_));
  OR4X1    g0535(.A(new_n1016_), .B(new_n985_), .C(new_n982_), .D(new_n932_), .Y(\V398(0) ));
  INVX1    g0536(.A(new_n920_), .Y(new_n1018_));
  INVX1    g0537(.A(\V16(0) ), .Y(new_n1019_));
  AND2X1   g0538(.A(\V15(0) ), .B(new_n1019_), .Y(new_n1020_));
  AND2X1   g0539(.A(\V15(0) ), .B(\V16(0) ), .Y(new_n1021_));
  NOR2X1   g0540(.A(new_n1021_), .B(new_n1020_), .Y(new_n1022_));
  AOI21X1  g0541(.A0(new_n996_), .A1(\V56(0) ), .B0(new_n1002_), .Y(new_n1023_));
  OAI21X1  g0542(.A0(new_n1009_), .A1(new_n1005_), .B0(new_n1023_), .Y(new_n1024_));
  NAND3X1  g0543(.A(new_n1024_), .B(new_n1022_), .C(new_n1018_), .Y(\V410(0) ));
  INVX1    g0544(.A(\V207(0) ), .Y(new_n1026_));
  AND2X1   g0545(.A(\V172(0) ), .B(\V56(0) ), .Y(new_n1027_));
  NOR2X1   g0546(.A(new_n1027_), .B(new_n1026_), .Y(new_n1028_));
  INVX1    g0547(.A(new_n1028_), .Y(new_n1029_));
  XOR2X1   g0548(.A(\V88(3) ), .B(new_n540_), .Y(new_n1030_));
  XOR2X1   g0549(.A(\V88(0) ), .B(\V88(1) ), .Y(new_n1031_));
  XOR2X1   g0550(.A(new_n1031_), .B(new_n1030_), .Y(new_n1032_));
  XOR2X1   g0551(.A(\V84(4) ), .B(\V84(5) ), .Y(new_n1033_));
  XOR2X1   g0552(.A(\V84(2) ), .B(\V84(3) ), .Y(new_n1034_));
  XOR2X1   g0553(.A(new_n1034_), .B(new_n1033_), .Y(new_n1035_));
  XOR2X1   g0554(.A(new_n1035_), .B(new_n1032_), .Y(new_n1036_));
  XOR2X1   g0555(.A(new_n1036_), .B(\V94(1) ), .Y(new_n1037_));
  XOR2X1   g0556(.A(\V84(0) ), .B(\V84(1) ), .Y(new_n1038_));
  XOR2X1   g0557(.A(\V78(4) ), .B(\V78(5) ), .Y(new_n1039_));
  XOR2X1   g0558(.A(new_n1039_), .B(new_n1038_), .Y(new_n1040_));
  INVX1    g0559(.A(\V78(2) ), .Y(new_n1041_));
  XOR2X1   g0560(.A(\V78(3) ), .B(new_n1041_), .Y(new_n1042_));
  XOR2X1   g0561(.A(\V78(0) ), .B(\V78(1) ), .Y(new_n1043_));
  XOR2X1   g0562(.A(new_n1043_), .B(new_n1042_), .Y(new_n1044_));
  XOR2X1   g0563(.A(new_n1044_), .B(new_n1040_), .Y(new_n1045_));
  XOR2X1   g0564(.A(new_n1045_), .B(\V94(0) ), .Y(new_n1046_));
  NAND3X1  g0565(.A(new_n485_), .B(new_n527_), .C(new_n501_), .Y(new_n1047_));
  NOR4X1   g0566(.A(new_n1047_), .B(new_n498_), .C(new_n496_), .D(new_n495_), .Y(new_n1048_));
  NOR4X1   g0567(.A(new_n499_), .B(new_n498_), .C(\V149(4) ), .D(\V149(6) ), .Y(new_n1049_));
  NOR3X1   g0568(.A(new_n1049_), .B(new_n1048_), .C(new_n529_), .Y(new_n1050_));
  INVX1    g0569(.A(new_n564_), .Y(new_n1051_));
  INVX1    g0570(.A(new_n536_), .Y(new_n1052_));
  NOR3X1   g0571(.A(new_n562_), .B(new_n1052_), .C(new_n1051_), .Y(new_n1053_));
  OAI22X1  g0572(.A0(new_n1053_), .A1(new_n493_), .B0(new_n1050_), .B1(new_n531_), .Y(new_n1054_));
  OAI21X1  g0573(.A0(new_n1046_), .A1(new_n1037_), .B0(new_n1054_), .Y(new_n1055_));
  INVX1    g0574(.A(new_n1022_), .Y(\V1757(0) ));
  XOR2X1   g0575(.A(new_n697_), .B(new_n704_), .Y(new_n1057_));
  XOR2X1   g0576(.A(new_n683_), .B(\V32(1) ), .Y(new_n1058_));
  NAND3X1  g0577(.A(new_n1058_), .B(new_n818_), .C(\V32(2) ), .Y(new_n1059_));
  NOR2X1   g0578(.A(new_n1059_), .B(new_n1057_), .Y(new_n1060_));
  AOI21X1  g0579(.A0(new_n697_), .A1(\V32(0) ), .B0(new_n1060_), .Y(new_n1061_));
  XOR2X1   g0580(.A(new_n644_), .B(\V32(2) ), .Y(new_n1062_));
  NOR4X1   g0581(.A(new_n1062_), .B(new_n1057_), .C(new_n626_), .D(new_n726_), .Y(new_n1063_));
  NOR3X1   g0582(.A(new_n1057_), .B(new_n832_), .C(new_n714_), .Y(new_n1064_));
  AOI21X1  g0583(.A0(new_n1063_), .A1(new_n1058_), .B0(new_n1064_), .Y(new_n1065_));
  OR4X1    g0584(.A(new_n493_), .B(new_n484_), .C(\V149(1) ), .D(\V149(0) ), .Y(new_n1066_));
  NOR4X1   g0585(.A(new_n499_), .B(new_n498_), .C(\V149(4) ), .D(new_n495_), .Y(new_n1067_));
  NOR2X1   g0586(.A(new_n500_), .B(\V174(0) ), .Y(new_n1068_));
  NOR4X1   g0587(.A(new_n502_), .B(new_n498_), .C(\V149(4) ), .D(new_n495_), .Y(new_n1069_));
  NOR4X1   g0588(.A(new_n1069_), .B(new_n1068_), .C(new_n1067_), .D(new_n1049_), .Y(new_n1070_));
  OAI21X1  g0589(.A0(new_n1070_), .A1(new_n531_), .B0(new_n1066_), .Y(new_n1071_));
  AOI21X1  g0590(.A0(new_n606_), .A1(new_n536_), .B0(new_n493_), .Y(new_n1072_));
  AND2X1   g0591(.A(new_n1072_), .B(new_n572_), .Y(new_n1073_));
  NOR3X1   g0592(.A(new_n510_), .B(\V292(0) ), .C(new_n991_), .Y(new_n1074_));
  NOR4X1   g0593(.A(new_n528_), .B(new_n498_), .C(\V149(4) ), .D(new_n495_), .Y(new_n1075_));
  AND2X1   g0594(.A(new_n1075_), .B(\V66(0) ), .Y(new_n1076_));
  NOR4X1   g0595(.A(new_n1076_), .B(new_n1074_), .C(new_n1073_), .D(new_n1071_), .Y(new_n1077_));
  AOI21X1  g0596(.A0(new_n1065_), .A1(new_n1061_), .B0(new_n1077_), .Y(new_n1078_));
  AND2X1   g0597(.A(\V66(0) ), .B(\V215(0) ), .Y(new_n1079_));
  OR4X1    g0598(.A(new_n1079_), .B(new_n578_), .C(\V214(0) ), .D(\V43(0) ), .Y(new_n1080_));
  NOR4X1   g0599(.A(new_n1080_), .B(new_n1078_), .C(\V1757(0) ), .D(new_n1014_), .Y(new_n1081_));
  NAND4X1  g0600(.A(new_n1081_), .B(new_n1055_), .C(new_n1029_), .D(\V423(0) ), .Y(new_n1082_));
  OR4X1    g0601(.A(new_n1082_), .B(new_n989_), .C(new_n987_), .D(new_n929_), .Y(new_n1083_));
  NOR4X1   g0602(.A(new_n1083_), .B(new_n985_), .C(new_n982_), .D(new_n932_), .Y(V432));
  AND2X1   g0603(.A(new_n529_), .B(\V62(0) ), .Y(new_n1085_));
  NOR3X1   g0604(.A(new_n562_), .B(new_n524_), .C(new_n486_), .Y(new_n1086_));
  NOR3X1   g0605(.A(new_n1086_), .B(new_n583_), .C(new_n493_), .Y(new_n1087_));
  INVX1    g0606(.A(new_n524_), .Y(new_n1088_));
  OAI21X1  g0607(.A0(new_n562_), .A1(new_n486_), .B0(\V241(0) ), .Y(new_n1089_));
  AND2X1   g0608(.A(new_n1089_), .B(new_n1088_), .Y(new_n1090_));
  NAND2X1  g0609(.A(new_n580_), .B(\V59(0) ), .Y(new_n1091_));
  OAI22X1  g0610(.A0(new_n1091_), .A1(new_n1090_), .B0(new_n530_), .B1(new_n531_), .Y(new_n1092_));
  NOR3X1   g0611(.A(new_n1092_), .B(new_n1087_), .C(\V270(0) ), .Y(new_n1093_));
  NOR3X1   g0612(.A(new_n1093_), .B(new_n1085_), .C(\V302(0) ), .Y(V630));
  OR2X1    g0613(.A(V630), .B(V432), .Y(\V435(0) ));
  INVX1    g0614(.A(\V14(0) ), .Y(new_n1096_));
  OR2X1    g0615(.A(new_n1096_), .B(\V271(0) ), .Y(\V500(0) ));
  INVX1    g0616(.A(new_n1067_), .Y(new_n1098_));
  NOR2X1   g0617(.A(new_n1069_), .B(new_n1067_), .Y(new_n1099_));
  OAI22X1  g0618(.A0(new_n1099_), .A1(new_n531_), .B0(new_n1098_), .B1(new_n1001_), .Y(new_n1100_));
  NAND2X1  g0619(.A(new_n537_), .B(\V59(0) ), .Y(new_n1101_));
  INVX1    g0620(.A(new_n559_), .Y(new_n1102_));
  OR2X1    g0621(.A(new_n1102_), .B(new_n486_), .Y(new_n1103_));
  NOR3X1   g0622(.A(new_n536_), .B(new_n538_), .C(new_n485_), .Y(new_n1104_));
  AND2X1   g0623(.A(new_n1055_), .B(new_n1049_), .Y(new_n1105_));
  NOR4X1   g0624(.A(new_n1105_), .B(new_n1104_), .C(new_n1103_), .D(new_n562_), .Y(new_n1106_));
  OAI21X1  g0625(.A0(new_n1106_), .A1(new_n531_), .B0(new_n1101_), .Y(new_n1107_));
  OR2X1    g0626(.A(new_n1107_), .B(new_n1100_), .Y(\V508(0) ));
  INVX1    g0627(.A(\V40(0) ), .Y(new_n1109_));
  INVX1    g0628(.A(\V45(0) ), .Y(new_n1110_));
  OAI21X1  g0629(.A0(new_n1110_), .A1(\V43(0) ), .B0(new_n1109_), .Y(\V511(0) ));
  XOR2X1   g0630(.A(\V44(0) ), .B(\V42(0) ), .Y(new_n1112_));
  XOR2X1   g0631(.A(\V38(0) ), .B(\V39(0) ), .Y(new_n1113_));
  NOR2X1   g0632(.A(new_n1113_), .B(new_n1112_), .Y(V512));
  NOR2X1   g0633(.A(new_n567_), .B(new_n1005_), .Y(new_n1115_));
  NOR3X1   g0634(.A(new_n994_), .B(new_n539_), .C(new_n1005_), .Y(new_n1116_));
  NOR3X1   g0635(.A(new_n994_), .B(new_n538_), .C(new_n531_), .Y(new_n1117_));
  AND2X1   g0636(.A(new_n993_), .B(\V56(0) ), .Y(new_n1118_));
  NOR3X1   g0637(.A(new_n554_), .B(new_n538_), .C(new_n1005_), .Y(new_n1119_));
  OR4X1    g0638(.A(new_n1119_), .B(new_n1118_), .C(new_n1117_), .D(new_n1002_), .Y(new_n1120_));
  NOR3X1   g0639(.A(new_n1120_), .B(new_n1116_), .C(new_n1115_), .Y(new_n1121_));
  INVX1    g0640(.A(\V214(0) ), .Y(\V1481(0) ));
  OAI21X1  g0641(.A0(new_n1027_), .A1(new_n1026_), .B0(\V1481(0) ), .Y(new_n1123_));
  NOR4X1   g0642(.A(new_n1123_), .B(new_n1121_), .C(new_n920_), .D(\V43(0) ), .Y(V527));
  NOR2X1   g0643(.A(new_n706_), .B(new_n606_), .Y(V537));
  AND2X1   g0644(.A(\V1213(1) ), .B(new_n562_), .Y(V538));
  NOR2X1   g0645(.A(new_n735_), .B(new_n606_), .Y(V539));
  NOR2X1   g0646(.A(new_n728_), .B(new_n606_), .Y(V540));
  INVX1    g0647(.A(\V257(6) ), .Y(new_n1129_));
  NOR4X1   g0648(.A(new_n588_), .B(new_n596_), .C(new_n595_), .D(new_n1129_), .Y(new_n1130_));
  NAND2X1  g0649(.A(new_n584_), .B(\V223(4) ), .Y(new_n1131_));
  NAND2X1  g0650(.A(new_n535_), .B(\V183(4) ), .Y(new_n1132_));
  MX2X1    g0651(.A(new_n1132_), .B(new_n1131_), .S0(new_n589_), .Y(new_n1133_));
  NOR4X1   g0652(.A(new_n1133_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1134_));
  OAI21X1  g0653(.A0(new_n1134_), .A1(new_n1130_), .B0(new_n575_), .Y(new_n1135_));
  NOR2X1   g0654(.A(new_n1135_), .B(new_n608_), .Y(new_n1136_));
  AND2X1   g0655(.A(new_n608_), .B(\V32(4) ), .Y(new_n1137_));
  MX2X1    g0656(.A(new_n1137_), .B(new_n1136_), .S0(new_n571_), .Y(\V1213(4) ));
  AND2X1   g0657(.A(\V1213(4) ), .B(new_n562_), .Y(V541));
  NAND2X1  g0658(.A(new_n578_), .B(\V257(0) ), .Y(new_n1140_));
  NOR3X1   g0659(.A(new_n1140_), .B(new_n588_), .C(new_n596_), .Y(new_n1141_));
  NAND2X1  g0660(.A(new_n584_), .B(\V223(5) ), .Y(new_n1142_));
  NAND2X1  g0661(.A(new_n535_), .B(\V183(5) ), .Y(new_n1143_));
  MX2X1    g0662(.A(new_n1143_), .B(new_n1142_), .S0(new_n589_), .Y(new_n1144_));
  NOR4X1   g0663(.A(new_n1144_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1145_));
  OAI21X1  g0664(.A0(new_n1145_), .A1(new_n1141_), .B0(new_n575_), .Y(new_n1146_));
  AND2X1   g0665(.A(new_n939_), .B(new_n574_), .Y(new_n1147_));
  INVX1    g0666(.A(new_n1147_), .Y(new_n1148_));
  AOI21X1  g0667(.A0(new_n1148_), .A1(new_n1146_), .B0(new_n608_), .Y(new_n1149_));
  AND2X1   g0668(.A(new_n608_), .B(\V32(5) ), .Y(new_n1150_));
  MX2X1    g0669(.A(new_n1150_), .B(new_n1149_), .S0(new_n571_), .Y(\V1213(5) ));
  AND2X1   g0670(.A(\V1213(5) ), .B(new_n562_), .Y(V542));
  NAND2X1  g0671(.A(new_n578_), .B(\V257(1) ), .Y(new_n1153_));
  NOR3X1   g0672(.A(new_n1153_), .B(new_n588_), .C(new_n596_), .Y(new_n1154_));
  NAND2X1  g0673(.A(new_n584_), .B(\V229(0) ), .Y(new_n1155_));
  NAND2X1  g0674(.A(new_n535_), .B(\V189(0) ), .Y(new_n1156_));
  MX2X1    g0675(.A(new_n1156_), .B(new_n1155_), .S0(new_n589_), .Y(new_n1157_));
  NOR4X1   g0676(.A(new_n1157_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1158_));
  OAI21X1  g0677(.A0(new_n1158_), .A1(new_n1154_), .B0(new_n575_), .Y(new_n1159_));
  AND2X1   g0678(.A(new_n602_), .B(new_n574_), .Y(new_n1160_));
  INVX1    g0679(.A(new_n1160_), .Y(new_n1161_));
  AOI21X1  g0680(.A0(new_n1161_), .A1(new_n1159_), .B0(new_n608_), .Y(new_n1162_));
  AND2X1   g0681(.A(new_n608_), .B(\V32(6) ), .Y(new_n1163_));
  MX2X1    g0682(.A(new_n1163_), .B(new_n1162_), .S0(new_n571_), .Y(\V1213(6) ));
  AND2X1   g0683(.A(\V1213(6) ), .B(new_n562_), .Y(V543));
  INVX1    g0684(.A(\V257(2) ), .Y(new_n1166_));
  NOR4X1   g0685(.A(new_n588_), .B(new_n596_), .C(new_n595_), .D(new_n1166_), .Y(new_n1167_));
  NAND2X1  g0686(.A(new_n584_), .B(\V229(1) ), .Y(new_n1168_));
  NAND2X1  g0687(.A(new_n535_), .B(\V189(1) ), .Y(new_n1169_));
  MX2X1    g0688(.A(new_n1169_), .B(new_n1168_), .S0(new_n589_), .Y(new_n1170_));
  NOR4X1   g0689(.A(new_n1170_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1171_));
  OAI21X1  g0690(.A0(new_n1171_), .A1(new_n1167_), .B0(new_n575_), .Y(new_n1172_));
  AOI21X1  g0691(.A0(new_n939_), .A1(new_n704_), .B0(new_n575_), .Y(new_n1173_));
  INVX1    g0692(.A(new_n1173_), .Y(new_n1174_));
  AOI21X1  g0693(.A0(new_n1174_), .A1(new_n1172_), .B0(new_n608_), .Y(new_n1175_));
  AND2X1   g0694(.A(new_n608_), .B(\V32(7) ), .Y(new_n1176_));
  MX2X1    g0695(.A(new_n1176_), .B(new_n1175_), .S0(new_n571_), .Y(\V1213(7) ));
  AND2X1   g0696(.A(\V1213(7) ), .B(new_n562_), .Y(V544));
  INVX1    g0697(.A(\V257(3) ), .Y(new_n1179_));
  NOR4X1   g0698(.A(new_n588_), .B(new_n596_), .C(new_n595_), .D(new_n1179_), .Y(new_n1180_));
  NAND2X1  g0699(.A(new_n584_), .B(\V229(2) ), .Y(new_n1181_));
  NAND2X1  g0700(.A(new_n535_), .B(\V189(2) ), .Y(new_n1182_));
  MX2X1    g0701(.A(new_n1182_), .B(new_n1181_), .S0(new_n589_), .Y(new_n1183_));
  NOR4X1   g0702(.A(new_n1183_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1184_));
  OAI21X1  g0703(.A0(new_n1184_), .A1(new_n1180_), .B0(new_n575_), .Y(new_n1185_));
  AOI21X1  g0704(.A0(new_n939_), .A1(new_n714_), .B0(new_n575_), .Y(new_n1186_));
  INVX1    g0705(.A(new_n1186_), .Y(new_n1187_));
  AOI21X1  g0706(.A0(new_n1187_), .A1(new_n1185_), .B0(new_n608_), .Y(new_n1188_));
  AND2X1   g0707(.A(new_n608_), .B(\V32(8) ), .Y(new_n1189_));
  MX2X1    g0708(.A(new_n1189_), .B(new_n1188_), .S0(new_n571_), .Y(\V1213(8) ));
  AND2X1   g0709(.A(\V1213(8) ), .B(new_n562_), .Y(V545));
  INVX1    g0710(.A(\V257(4) ), .Y(new_n1192_));
  NOR4X1   g0711(.A(new_n588_), .B(new_n596_), .C(new_n595_), .D(new_n1192_), .Y(new_n1193_));
  NAND2X1  g0712(.A(new_n584_), .B(\V229(3) ), .Y(new_n1194_));
  NAND2X1  g0713(.A(new_n535_), .B(\V189(3) ), .Y(new_n1195_));
  MX2X1    g0714(.A(new_n1195_), .B(new_n1194_), .S0(new_n589_), .Y(new_n1196_));
  NOR4X1   g0715(.A(new_n1196_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1197_));
  OAI21X1  g0716(.A0(new_n1197_), .A1(new_n1193_), .B0(new_n575_), .Y(new_n1198_));
  AOI21X1  g0717(.A0(new_n939_), .A1(new_n733_), .B0(new_n575_), .Y(new_n1199_));
  INVX1    g0718(.A(new_n1199_), .Y(new_n1200_));
  AOI21X1  g0719(.A0(new_n1200_), .A1(new_n1198_), .B0(new_n608_), .Y(new_n1201_));
  AND2X1   g0720(.A(new_n608_), .B(\V32(9) ), .Y(new_n1202_));
  MX2X1    g0721(.A(new_n1202_), .B(new_n1201_), .S0(new_n571_), .Y(\V1213(9) ));
  AND2X1   g0722(.A(\V1213(9) ), .B(new_n562_), .Y(V546));
  NAND2X1  g0723(.A(new_n578_), .B(\V257(5) ), .Y(new_n1205_));
  NOR3X1   g0724(.A(new_n1205_), .B(new_n588_), .C(new_n596_), .Y(new_n1206_));
  NAND2X1  g0725(.A(new_n584_), .B(\V229(4) ), .Y(new_n1207_));
  NAND2X1  g0726(.A(new_n535_), .B(\V189(4) ), .Y(new_n1208_));
  MX2X1    g0727(.A(new_n1208_), .B(new_n1207_), .S0(new_n589_), .Y(new_n1209_));
  NOR4X1   g0728(.A(new_n1209_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1210_));
  OAI21X1  g0729(.A0(new_n1210_), .A1(new_n1206_), .B0(new_n575_), .Y(new_n1211_));
  MX2X1    g0730(.A(\V32(3) ), .B(\V32(0) ), .S0(new_n602_), .Y(new_n1212_));
  AND2X1   g0731(.A(new_n1212_), .B(new_n574_), .Y(new_n1213_));
  INVX1    g0732(.A(new_n1213_), .Y(new_n1214_));
  AOI21X1  g0733(.A0(new_n1214_), .A1(new_n1211_), .B0(new_n608_), .Y(new_n1215_));
  AND2X1   g0734(.A(new_n608_), .B(\V32(10) ), .Y(new_n1216_));
  MX2X1    g0735(.A(new_n1216_), .B(new_n1215_), .S0(new_n571_), .Y(\V1213(10) ));
  AND2X1   g0736(.A(\V1213(10) ), .B(new_n562_), .Y(V547));
  NAND2X1  g0737(.A(new_n584_), .B(\V229(5) ), .Y(new_n1219_));
  NAND2X1  g0738(.A(new_n535_), .B(\V189(5) ), .Y(new_n1220_));
  MX2X1    g0739(.A(new_n1220_), .B(new_n1219_), .S0(new_n589_), .Y(new_n1221_));
  NOR4X1   g0740(.A(new_n1221_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1222_));
  OAI21X1  g0741(.A0(new_n1222_), .A1(new_n1130_), .B0(new_n575_), .Y(new_n1223_));
  MX2X1    g0742(.A(\V32(4) ), .B(\V32(1) ), .S0(new_n602_), .Y(new_n1224_));
  AND2X1   g0743(.A(new_n1224_), .B(new_n574_), .Y(new_n1225_));
  INVX1    g0744(.A(new_n1225_), .Y(new_n1226_));
  AOI21X1  g0745(.A0(new_n1226_), .A1(new_n1223_), .B0(new_n608_), .Y(new_n1227_));
  AND2X1   g0746(.A(new_n608_), .B(\V32(11) ), .Y(new_n1228_));
  MX2X1    g0747(.A(new_n1228_), .B(new_n1227_), .S0(new_n571_), .Y(\V1213(11) ));
  AND2X1   g0748(.A(\V1213(11) ), .B(new_n562_), .Y(V548));
  AND2X1   g0749(.A(\V802(0) ), .B(new_n486_), .Y(new_n1231_));
  NOR3X1   g0750(.A(new_n589_), .B(new_n580_), .C(\V802(0) ), .Y(new_n1232_));
  INVX1    g0751(.A(\V134(1) ), .Y(new_n1233_));
  NAND4X1  g0752(.A(new_n927_), .B(\V194(0) ), .C(\V199(1) ), .D(\V199(3) ), .Y(new_n1234_));
  INVX1    g0753(.A(\V271(0) ), .Y(new_n1235_));
  NOR3X1   g0754(.A(new_n529_), .B(\V274(0) ), .C(new_n1235_), .Y(new_n1236_));
  NAND4X1  g0755(.A(new_n1236_), .B(new_n1234_), .C(new_n580_), .D(\V134(0) ), .Y(new_n1237_));
  NOR2X1   g0756(.A(new_n1237_), .B(new_n1233_), .Y(new_n1238_));
  NOR2X1   g0757(.A(new_n1238_), .B(new_n1232_), .Y(new_n1239_));
  NAND4X1  g0758(.A(new_n1239_), .B(\V1243(9) ), .C(new_n562_), .D(\V802(0) ), .Y(new_n1240_));
  NOR4X1   g0759(.A(new_n506_), .B(new_n493_), .C(\V149(3) ), .D(\V174(0) ), .Y(new_n1241_));
  OR4X1    g0760(.A(new_n1241_), .B(new_n1239_), .C(new_n1231_), .D(\V199(4) ), .Y(new_n1242_));
  OAI21X1  g0761(.A0(new_n1240_), .A1(new_n1231_), .B0(new_n1242_), .Y(\V572(9) ));
  NAND4X1  g0762(.A(new_n1239_), .B(\V1243(8) ), .C(new_n562_), .D(\V802(0) ), .Y(new_n1244_));
  INVX1    g0763(.A(\V199(3) ), .Y(new_n1245_));
  XOR2X1   g0764(.A(new_n1245_), .B(\V199(4) ), .Y(new_n1246_));
  OR4X1    g0765(.A(new_n1246_), .B(new_n1241_), .C(new_n1239_), .D(new_n1231_), .Y(new_n1247_));
  OAI21X1  g0766(.A0(new_n1244_), .A1(new_n1231_), .B0(new_n1247_), .Y(\V572(8) ));
  NAND4X1  g0767(.A(new_n1239_), .B(\V1243(7) ), .C(new_n562_), .D(\V802(0) ), .Y(new_n1249_));
  NAND2X1  g0768(.A(\V199(3) ), .B(\V199(4) ), .Y(new_n1250_));
  XOR2X1   g0769(.A(new_n1250_), .B(\V199(2) ), .Y(new_n1251_));
  OR4X1    g0770(.A(new_n1251_), .B(new_n1241_), .C(new_n1239_), .D(new_n1231_), .Y(new_n1252_));
  OAI21X1  g0771(.A0(new_n1249_), .A1(new_n1231_), .B0(new_n1252_), .Y(\V572(7) ));
  NAND2X1  g0772(.A(new_n584_), .B(\V239(1) ), .Y(new_n1254_));
  NAND2X1  g0773(.A(new_n535_), .B(\V199(1) ), .Y(new_n1255_));
  MX2X1    g0774(.A(new_n1255_), .B(new_n1254_), .S0(new_n589_), .Y(new_n1256_));
  OR4X1    g0775(.A(new_n1256_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1257_));
  INVX1    g0776(.A(\V32(8) ), .Y(new_n1258_));
  MX2X1    g0777(.A(new_n938_), .B(new_n1258_), .S0(new_n602_), .Y(new_n1259_));
  MX2X1    g0778(.A(new_n1259_), .B(new_n1257_), .S0(new_n575_), .Y(new_n1260_));
  NOR2X1   g0779(.A(new_n1260_), .B(new_n608_), .Y(new_n1261_));
  AND2X1   g0780(.A(new_n608_), .B(\V84(4) ), .Y(new_n1262_));
  MX2X1    g0781(.A(new_n1262_), .B(new_n1261_), .S0(new_n571_), .Y(\V1243(6) ));
  NAND4X1  g0782(.A(\V1243(6) ), .B(new_n1239_), .C(new_n562_), .D(\V802(0) ), .Y(new_n1264_));
  NAND3X1  g0783(.A(\V199(2) ), .B(\V199(3) ), .C(\V199(4) ), .Y(new_n1265_));
  XOR2X1   g0784(.A(new_n1265_), .B(\V199(1) ), .Y(new_n1266_));
  OR4X1    g0785(.A(new_n1266_), .B(new_n1241_), .C(new_n1239_), .D(new_n1231_), .Y(new_n1267_));
  OAI21X1  g0786(.A0(new_n1264_), .A1(new_n1231_), .B0(new_n1267_), .Y(\V572(6) ));
  NAND2X1  g0787(.A(new_n584_), .B(\V239(0) ), .Y(new_n1269_));
  NAND2X1  g0788(.A(new_n535_), .B(\V199(0) ), .Y(new_n1270_));
  MX2X1    g0789(.A(new_n1270_), .B(new_n1269_), .S0(new_n589_), .Y(new_n1271_));
  OR4X1    g0790(.A(new_n1271_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1272_));
  INVX1    g0791(.A(\V32(7) ), .Y(new_n1273_));
  MX2X1    g0792(.A(new_n961_), .B(new_n1273_), .S0(new_n602_), .Y(new_n1274_));
  MX2X1    g0793(.A(new_n1274_), .B(new_n1272_), .S0(new_n575_), .Y(new_n1275_));
  NOR2X1   g0794(.A(new_n1275_), .B(new_n608_), .Y(new_n1276_));
  AND2X1   g0795(.A(new_n608_), .B(\V84(3) ), .Y(new_n1277_));
  MX2X1    g0796(.A(new_n1277_), .B(new_n1276_), .S0(new_n571_), .Y(\V1243(5) ));
  NAND4X1  g0797(.A(\V1243(5) ), .B(new_n1239_), .C(new_n562_), .D(\V802(0) ), .Y(new_n1279_));
  NAND4X1  g0798(.A(\V199(1) ), .B(\V199(2) ), .C(\V199(3) ), .D(\V199(4) ), .Y(new_n1280_));
  XOR2X1   g0799(.A(new_n1280_), .B(\V199(0) ), .Y(new_n1281_));
  OR4X1    g0800(.A(new_n1281_), .B(new_n1241_), .C(new_n1239_), .D(new_n1231_), .Y(new_n1282_));
  OAI21X1  g0801(.A0(new_n1279_), .A1(new_n1231_), .B0(new_n1282_), .Y(\V572(5) ));
  NAND2X1  g0802(.A(new_n584_), .B(\V234(4) ), .Y(new_n1284_));
  NAND2X1  g0803(.A(new_n535_), .B(\V194(4) ), .Y(new_n1285_));
  MX2X1    g0804(.A(new_n1285_), .B(new_n1284_), .S0(new_n589_), .Y(new_n1286_));
  OR4X1    g0805(.A(new_n1286_), .B(new_n588_), .C(new_n587_), .D(new_n578_), .Y(new_n1287_));
  INVX1    g0806(.A(\V32(6) ), .Y(new_n1288_));
  MX2X1    g0807(.A(new_n950_), .B(new_n1288_), .S0(new_n602_), .Y(new_n1289_));
  MX2X1    g0808(.A(new_n1289_), .B(new_n1287_), .S0(new_n575_), .Y(new_n1290_));
  NOR2X1   g0809(.A(new_n1290_), .B(new_n608_), .Y(new_n1291_));
  AND2X1   g0810(.A(new_n608_), .B(\V84(2) ), .Y(new_n1292_));
  MX2X1    g0811(.A(new_n1292_), .B(new_n1291_), .S0(new_n571_), .Y(\V1243(4) ));
  NAND4X1  g0812(.A(\V1243(4) ), .B(new_n1239_), .C(new_n562_), .D(\V802(0) ), .Y(new_n1294_));
  INVX1    g0813(.A(\V199(1) ), .Y(new_n1295_));
  NAND3X1  g0814(.A(\V199(0) ), .B(\V199(2) ), .C(\V199(4) ), .Y(new_n1296_));
  NOR3X1   g0815(.A(new_n1296_), .B(new_n1295_), .C(new_n1245_), .Y(new_n1297_));
  XOR2X1   g0816(.A(new_n1297_), .B(new_n923_), .Y(new_n1298_));
  OR4X1    g0817(.A(new_n1298_), .B(new_n1241_), .C(new_n1239_), .D(new_n1231_), .Y(new_n1299_));
  OAI21X1  g0818(.A0(new_n1294_), .A1(new_n1231_), .B0(new_n1299_), .Y(\V572(4) ));
  INVX1    g0819(.A(new_n1239_), .Y(new_n1301_));
  INVX1    g0820(.A(new_n577_), .Y(new_n1302_));
  NAND2X1  g0821(.A(new_n584_), .B(\V234(3) ), .Y(new_n1303_));
  NAND2X1  g0822(.A(new_n535_), .B(\V194(3) ), .Y(new_n1304_));
  MX2X1    g0823(.A(new_n1304_), .B(new_n1303_), .S0(new_n589_), .Y(new_n1305_));
  OR4X1    g0824(.A(new_n1305_), .B(new_n588_), .C(new_n1302_), .D(\V262(0) ), .Y(new_n1306_));
  NOR4X1   g0825(.A(new_n580_), .B(new_n579_), .C(new_n501_), .D(\V59(0) ), .Y(new_n1307_));
  NAND4X1  g0826(.A(new_n1307_), .B(new_n587_), .C(new_n577_), .D(new_n576_), .Y(new_n1308_));
  OAI21X1  g0827(.A0(new_n1306_), .A1(new_n587_), .B0(new_n1308_), .Y(new_n1309_));
  MX2X1    g0828(.A(\V32(8) ), .B(\V32(5) ), .S0(new_n602_), .Y(new_n1310_));
  MX2X1    g0829(.A(new_n1310_), .B(new_n1309_), .S0(new_n575_), .Y(new_n1311_));
  OAI21X1  g0830(.A0(new_n607_), .A1(new_n571_), .B0(new_n1311_), .Y(new_n1312_));
  AND2X1   g0831(.A(new_n608_), .B(\V84(1) ), .Y(new_n1313_));
  INVX1    g0832(.A(new_n1313_), .Y(new_n1314_));
  MX2X1    g0833(.A(new_n1314_), .B(new_n1312_), .S0(new_n571_), .Y(new_n1315_));
  OR4X1    g0834(.A(new_n1315_), .B(new_n1301_), .C(new_n606_), .D(new_n493_), .Y(new_n1316_));
  NOR4X1   g0835(.A(new_n1301_), .B(new_n493_), .C(new_n579_), .D(new_n501_), .Y(new_n1317_));
  OR4X1    g0836(.A(new_n1296_), .B(new_n923_), .C(new_n1295_), .D(new_n1245_), .Y(new_n1318_));
  XOR2X1   g0837(.A(new_n1318_), .B(\V194(3) ), .Y(new_n1319_));
  NOR3X1   g0838(.A(new_n1319_), .B(new_n1239_), .C(new_n1231_), .Y(new_n1320_));
  OAI22X1  g0839(.A0(new_n1320_), .A1(new_n1317_), .B0(new_n606_), .B1(new_n493_), .Y(new_n1321_));
  OAI21X1  g0840(.A0(new_n1316_), .A1(new_n1231_), .B0(new_n1321_), .Y(\V572(3) ));
  NAND2X1  g0841(.A(new_n584_), .B(\V234(2) ), .Y(new_n1323_));
  NAND2X1  g0842(.A(new_n535_), .B(\V194(2) ), .Y(new_n1324_));
  MX2X1    g0843(.A(new_n1324_), .B(new_n1323_), .S0(new_n589_), .Y(new_n1325_));
  OR4X1    g0844(.A(new_n1325_), .B(new_n588_), .C(new_n1302_), .D(\V262(0) ), .Y(new_n1326_));
  NOR4X1   g0845(.A(new_n580_), .B(new_n579_), .C(new_n495_), .D(\V59(0) ), .Y(new_n1327_));
  NAND4X1  g0846(.A(new_n1327_), .B(new_n587_), .C(new_n577_), .D(new_n576_), .Y(new_n1328_));
  OAI21X1  g0847(.A0(new_n1326_), .A1(new_n587_), .B0(new_n1328_), .Y(new_n1329_));
  MX2X1    g0848(.A(\V32(7) ), .B(\V32(4) ), .S0(new_n602_), .Y(new_n1330_));
  MX2X1    g0849(.A(new_n1330_), .B(new_n1329_), .S0(new_n575_), .Y(new_n1331_));
  OAI21X1  g0850(.A0(new_n607_), .A1(new_n571_), .B0(new_n1331_), .Y(new_n1332_));
  AND2X1   g0851(.A(new_n608_), .B(\V84(0) ), .Y(new_n1333_));
  INVX1    g0852(.A(new_n1333_), .Y(new_n1334_));
  MX2X1    g0853(.A(new_n1334_), .B(new_n1332_), .S0(new_n571_), .Y(new_n1335_));
  OR4X1    g0854(.A(new_n1335_), .B(new_n1301_), .C(new_n606_), .D(new_n493_), .Y(new_n1336_));
  NOR4X1   g0855(.A(new_n1301_), .B(new_n493_), .C(new_n579_), .D(new_n495_), .Y(new_n1337_));
  NOR4X1   g0856(.A(new_n926_), .B(new_n923_), .C(new_n1295_), .D(new_n1245_), .Y(new_n1338_));
  XOR2X1   g0857(.A(new_n1338_), .B(new_n924_), .Y(new_n1339_));
  NOR3X1   g0858(.A(new_n1339_), .B(new_n1239_), .C(new_n1231_), .Y(new_n1340_));
  OAI22X1  g0859(.A0(new_n1340_), .A1(new_n1337_), .B0(new_n606_), .B1(new_n493_), .Y(new_n1341_));
  OAI21X1  g0860(.A0(new_n1336_), .A1(new_n1231_), .B0(new_n1341_), .Y(\V572(2) ));
  NAND2X1  g0861(.A(new_n584_), .B(\V234(1) ), .Y(new_n1343_));
  NAND2X1  g0862(.A(new_n535_), .B(\V194(1) ), .Y(new_n1344_));
  MX2X1    g0863(.A(new_n1344_), .B(new_n1343_), .S0(new_n589_), .Y(new_n1345_));
  OR4X1    g0864(.A(new_n1345_), .B(new_n588_), .C(new_n1302_), .D(\V262(0) ), .Y(new_n1346_));
  NOR4X1   g0865(.A(new_n580_), .B(new_n579_), .C(new_n527_), .D(\V59(0) ), .Y(new_n1347_));
  NAND4X1  g0866(.A(new_n1347_), .B(new_n587_), .C(new_n577_), .D(new_n576_), .Y(new_n1348_));
  OAI21X1  g0867(.A0(new_n1346_), .A1(new_n587_), .B0(new_n1348_), .Y(new_n1349_));
  MX2X1    g0868(.A(\V32(6) ), .B(\V32(3) ), .S0(new_n602_), .Y(new_n1350_));
  MX2X1    g0869(.A(new_n1350_), .B(new_n1349_), .S0(new_n575_), .Y(new_n1351_));
  OAI21X1  g0870(.A0(new_n607_), .A1(new_n571_), .B0(new_n1351_), .Y(new_n1352_));
  AND2X1   g0871(.A(new_n608_), .B(\V78(5) ), .Y(new_n1353_));
  INVX1    g0872(.A(new_n1353_), .Y(new_n1354_));
  MX2X1    g0873(.A(new_n1354_), .B(new_n1352_), .S0(new_n571_), .Y(new_n1355_));
  OR4X1    g0874(.A(new_n1355_), .B(new_n1301_), .C(new_n606_), .D(new_n493_), .Y(new_n1356_));
  NOR4X1   g0875(.A(new_n1301_), .B(new_n493_), .C(new_n579_), .D(new_n527_), .Y(new_n1357_));
  NOR4X1   g0876(.A(new_n926_), .B(new_n924_), .C(new_n923_), .D(new_n1295_), .Y(new_n1358_));
  AND2X1   g0877(.A(new_n1358_), .B(\V199(3) ), .Y(new_n1359_));
  XOR2X1   g0878(.A(new_n1359_), .B(new_n925_), .Y(new_n1360_));
  NOR3X1   g0879(.A(new_n1360_), .B(new_n1239_), .C(new_n1231_), .Y(new_n1361_));
  OAI22X1  g0880(.A0(new_n1361_), .A1(new_n1357_), .B0(new_n606_), .B1(new_n493_), .Y(new_n1362_));
  OAI21X1  g0881(.A0(new_n1356_), .A1(new_n1231_), .B0(new_n1362_), .Y(\V572(1) ));
  NAND4X1  g0882(.A(new_n1239_), .B(\V1243(0) ), .C(new_n562_), .D(\V802(0) ), .Y(new_n1364_));
  NOR4X1   g0883(.A(new_n1301_), .B(new_n493_), .C(new_n579_), .D(new_n496_), .Y(new_n1365_));
  XOR2X1   g0884(.A(new_n928_), .B(\V194(0) ), .Y(new_n1366_));
  NOR3X1   g0885(.A(new_n1366_), .B(new_n1239_), .C(new_n1231_), .Y(new_n1367_));
  OAI22X1  g0886(.A0(new_n1367_), .A1(new_n1365_), .B0(new_n606_), .B1(new_n493_), .Y(new_n1368_));
  OAI21X1  g0887(.A0(new_n1364_), .A1(new_n1231_), .B0(new_n1368_), .Y(\V572(0) ));
  INVX1    g0888(.A(\V34(0) ), .Y(\V585(0) ));
  INVX1    g0889(.A(new_n589_), .Y(new_n1371_));
  AOI21X1  g0890(.A0(new_n1371_), .A1(\V802(0) ), .B0(\V243(0) ), .Y(V587));
  INVX1    g0891(.A(\V244(0) ), .Y(new_n1373_));
  OR2X1    g0892(.A(new_n1373_), .B(\V243(0) ), .Y(new_n1374_));
  INVX1    g0893(.A(\V243(0) ), .Y(new_n1375_));
  OR2X1    g0894(.A(\V244(0) ), .B(new_n1375_), .Y(new_n1376_));
  AOI22X1  g0895(.A0(new_n1376_), .A1(new_n1374_), .B0(new_n1371_), .B1(\V802(0) ), .Y(\V591(0) ));
  OAI21X1  g0896(.A0(new_n1373_), .A1(new_n1375_), .B0(\V245(0) ), .Y(new_n1378_));
  NAND2X1  g0897(.A(\V244(0) ), .B(\V243(0) ), .Y(new_n1379_));
  OR2X1    g0898(.A(new_n1379_), .B(\V245(0) ), .Y(new_n1380_));
  AOI22X1  g0899(.A0(new_n1380_), .A1(new_n1378_), .B0(new_n1371_), .B1(\V802(0) ), .Y(\V597(0) ));
  NAND3X1  g0900(.A(\V245(0) ), .B(\V244(0) ), .C(\V243(0) ), .Y(new_n1382_));
  NAND2X1  g0901(.A(new_n1382_), .B(\V246(0) ), .Y(new_n1383_));
  OR2X1    g0902(.A(new_n1382_), .B(\V246(0) ), .Y(new_n1384_));
  AOI22X1  g0903(.A0(new_n1384_), .A1(new_n1383_), .B0(new_n1371_), .B1(\V802(0) ), .Y(\V603(0) ));
  NAND2X1  g0904(.A(new_n931_), .B(\V247(0) ), .Y(new_n1386_));
  OR2X1    g0905(.A(new_n931_), .B(\V247(0) ), .Y(new_n1387_));
  AOI22X1  g0906(.A0(new_n1387_), .A1(new_n1386_), .B0(new_n1371_), .B1(\V802(0) ), .Y(\V609(0) ));
  AOI21X1  g0907(.A0(new_n1055_), .A1(new_n1049_), .B0(new_n537_), .Y(new_n1389_));
  NOR4X1   g0908(.A(new_n1389_), .B(new_n920_), .C(\V214(0) ), .D(new_n1005_), .Y(new_n1390_));
  NOR4X1   g0909(.A(new_n1098_), .B(new_n920_), .C(\V214(0) ), .D(new_n1001_), .Y(new_n1391_));
  OR2X1    g0910(.A(new_n1028_), .B(new_n920_), .Y(new_n1392_));
  NOR4X1   g0911(.A(new_n1392_), .B(new_n1106_), .C(\V214(0) ), .D(new_n531_), .Y(new_n1393_));
  NOR3X1   g0912(.A(new_n1393_), .B(new_n1391_), .C(new_n1390_), .Y(V620));
  INVX1    g0913(.A(\V293(0) ), .Y(new_n1395_));
  XOR2X1   g0914(.A(\V41(0) ), .B(\V45(0) ), .Y(new_n1396_));
  NOR2X1   g0915(.A(new_n1396_), .B(new_n1395_), .Y(V621));
  NAND3X1  g0916(.A(\V202(0) ), .B(\V274(0) ), .C(new_n1235_), .Y(new_n1398_));
  NAND2X1  g0917(.A(\V269(0) ), .B(\V271(0) ), .Y(new_n1399_));
  AND2X1   g0918(.A(new_n1399_), .B(new_n1398_), .Y(\V634(0) ));
  INVX1    g0919(.A(\V274(0) ), .Y(new_n1401_));
  OAI21X1  g0920(.A0(\V202(0) ), .A1(new_n1401_), .B0(new_n1235_), .Y(\V640(0) ));
  INVX1    g0921(.A(new_n541_), .Y(V707));
  INVX1    g0922(.A(new_n572_), .Y(V763));
  NOR4X1   g0923(.A(new_n1090_), .B(new_n580_), .C(\V802(0) ), .D(\V1833(0) ), .Y(new_n1405_));
  INVX1    g0924(.A(\V272(0) ), .Y(new_n1406_));
  NAND4X1  g0925(.A(new_n493_), .B(\V134(0) ), .C(\V134(1) ), .D(\V242(0) ), .Y(new_n1407_));
  NOR4X1   g0926(.A(new_n1407_), .B(new_n583_), .C(new_n1406_), .D(\V275(0) ), .Y(new_n1408_));
  INVX1    g0927(.A(\V242(0) ), .Y(new_n1409_));
  NOR2X1   g0928(.A(new_n562_), .B(new_n486_), .Y(new_n1410_));
  OAI21X1  g0929(.A0(new_n1410_), .A1(new_n531_), .B0(new_n583_), .Y(new_n1411_));
  NOR4X1   g0930(.A(new_n1411_), .B(new_n589_), .C(\V802(0) ), .D(new_n1409_), .Y(new_n1412_));
  OR4X1    g0931(.A(new_n1090_), .B(\V802(0) ), .C(new_n1406_), .D(\V1833(0) ), .Y(new_n1413_));
  OR2X1    g0932(.A(new_n1413_), .B(\V275(0) ), .Y(new_n1414_));
  INVX1    g0933(.A(new_n1068_), .Y(new_n1415_));
  NOR4X1   g0934(.A(new_n1415_), .B(new_n1029_), .C(new_n1051_), .D(new_n1005_), .Y(new_n1416_));
  INVX1    g0935(.A(\V67(0) ), .Y(new_n1417_));
  INVX1    g0936(.A(\V172(0) ), .Y(new_n1418_));
  NOR3X1   g0937(.A(new_n1418_), .B(new_n1417_), .C(new_n990_), .Y(new_n1419_));
  NOR4X1   g0938(.A(new_n502_), .B(new_n498_), .C(\V149(4) ), .D(\V149(6) ), .Y(new_n1420_));
  NAND2X1  g0939(.A(new_n1028_), .B(new_n564_), .Y(new_n1421_));
  NOR4X1   g0940(.A(new_n1421_), .B(new_n1420_), .C(new_n1068_), .D(new_n538_), .Y(new_n1422_));
  NAND4X1  g0941(.A(new_n1420_), .B(new_n1028_), .C(new_n564_), .D(\V62(0) ), .Y(new_n1423_));
  NAND4X1  g0942(.A(new_n1028_), .B(new_n538_), .C(new_n564_), .D(\V59(0) ), .Y(new_n1424_));
  NAND3X1  g0943(.A(new_n1424_), .B(new_n1423_), .C(\V1481(0) ), .Y(new_n1425_));
  NOR4X1   g0944(.A(new_n1425_), .B(new_n1422_), .C(new_n1419_), .D(new_n1416_), .Y(new_n1426_));
  OAI21X1  g0945(.A0(new_n1414_), .A1(new_n583_), .B0(new_n1426_), .Y(new_n1427_));
  NOR4X1   g0946(.A(new_n1427_), .B(new_n1412_), .C(new_n1408_), .D(new_n1405_), .Y(new_n1428_));
  INVX1    g0947(.A(new_n1428_), .Y(new_n1429_));
  INVX1    g0948(.A(\V165(7) ), .Y(new_n1430_));
  NOR3X1   g0949(.A(new_n1018_), .B(\V290(0) ), .C(new_n1430_), .Y(new_n1431_));
  NOR4X1   g0950(.A(new_n1431_), .B(new_n1429_), .C(new_n988_), .D(\V302(0) ), .Y(new_n1432_));
  NAND4X1  g0951(.A(new_n1432_), .B(new_n1302_), .C(V763), .D(\V70(0) ), .Y(new_n1433_));
  NOR2X1   g0952(.A(new_n1433_), .B(new_n1096_), .Y(V775));
  INVX1    g0953(.A(\V10(0) ), .Y(new_n1435_));
  INVX1    g0954(.A(\V6(0) ), .Y(new_n1436_));
  NOR3X1   g0955(.A(new_n1436_), .B(\V13(0) ), .C(new_n1435_), .Y(V779));
  INVX1    g0956(.A(\V12(0) ), .Y(new_n1438_));
  INVX1    g0957(.A(\V174(0) ), .Y(new_n1439_));
  AOI21X1  g0958(.A0(new_n503_), .A1(new_n500_), .B0(new_n531_), .Y(new_n1440_));
  AOI21X1  g0959(.A0(new_n1440_), .A1(new_n1439_), .B0(\V52(0) ), .Y(new_n1441_));
  NOR3X1   g0960(.A(new_n1441_), .B(new_n1438_), .C(new_n1436_), .Y(V781));
  INVX1    g0961(.A(\V7(0) ), .Y(new_n1443_));
  NOR3X1   g0962(.A(new_n1443_), .B(\V13(0) ), .C(new_n1435_), .Y(V782));
  AND2X1   g0963(.A(\V11(0) ), .B(\V5(0) ), .Y(V783));
  AND2X1   g0964(.A(\V11(0) ), .B(\V7(0) ), .Y(V784));
  INVX1    g0965(.A(\V9(0) ), .Y(new_n1447_));
  INVX1    g0966(.A(\V4(0) ), .Y(new_n1448_));
  NOR3X1   g0967(.A(new_n912_), .B(new_n1448_), .C(new_n1447_), .Y(V789));
  AND2X1   g0968(.A(new_n1422_), .B(new_n1018_), .Y(new_n1450_));
  AND2X1   g0969(.A(new_n1416_), .B(new_n1018_), .Y(new_n1451_));
  INVX1    g0970(.A(\V290(0) ), .Y(new_n1452_));
  NOR4X1   g0971(.A(new_n1452_), .B(new_n513_), .C(\V165(2) ), .D(new_n511_), .Y(new_n1453_));
  OAI21X1  g0972(.A0(new_n1424_), .A1(new_n920_), .B0(new_n1423_), .Y(new_n1454_));
  NOR4X1   g0973(.A(new_n1454_), .B(new_n1453_), .C(new_n1451_), .D(new_n1450_), .Y(new_n1455_));
  INVX1    g0974(.A(new_n1455_), .Y(\V1741(0) ));
  OR2X1    g0975(.A(new_n1069_), .B(new_n1049_), .Y(new_n1457_));
  NOR4X1   g0976(.A(new_n528_), .B(new_n498_), .C(\V149(4) ), .D(\V149(6) ), .Y(new_n1458_));
  NOR4X1   g0977(.A(new_n528_), .B(new_n498_), .C(new_n496_), .D(\V149(6) ), .Y(new_n1459_));
  NOR4X1   g0978(.A(new_n1047_), .B(new_n498_), .C(\V149(4) ), .D(new_n495_), .Y(new_n1460_));
  INVX1    g0979(.A(\V258(0) ), .Y(new_n1461_));
  OR4X1    g0980(.A(new_n595_), .B(\V260(0) ), .C(\V259(0) ), .D(\V59(0) ), .Y(new_n1462_));
  NOR4X1   g0981(.A(new_n1047_), .B(new_n498_), .C(new_n496_), .D(\V149(6) ), .Y(new_n1463_));
  NOR4X1   g0982(.A(new_n499_), .B(new_n498_), .C(new_n496_), .D(\V149(6) ), .Y(new_n1464_));
  NOR3X1   g0983(.A(new_n1464_), .B(new_n1463_), .C(new_n1048_), .Y(new_n1465_));
  OAI21X1  g0984(.A0(new_n1462_), .A1(new_n1461_), .B0(new_n1465_), .Y(new_n1466_));
  NOR4X1   g0985(.A(new_n1466_), .B(new_n1460_), .C(new_n1459_), .D(new_n1458_), .Y(new_n1467_));
  NAND2X1  g0986(.A(new_n1067_), .B(\V65(0) ), .Y(new_n1468_));
  OAI21X1  g0987(.A0(new_n1467_), .A1(new_n531_), .B0(new_n1468_), .Y(new_n1469_));
  AOI21X1  g0988(.A0(new_n1457_), .A1(\V62(0) ), .B0(new_n1469_), .Y(new_n1470_));
  NOR3X1   g0989(.A(new_n1470_), .B(\V1741(0) ), .C(new_n988_), .Y(new_n1471_));
  NOR2X1   g0990(.A(new_n920_), .B(new_n1452_), .Y(new_n1472_));
  OR4X1    g0991(.A(new_n1472_), .B(new_n1471_), .C(\V302(0) ), .D(\V289(0) ), .Y(new_n1473_));
  INVX1    g0992(.A(new_n1090_), .Y(new_n1474_));
  INVX1    g0993(.A(new_n1432_), .Y(new_n1475_));
  OAI21X1  g0994(.A0(new_n1475_), .A1(new_n916_), .B0(new_n1474_), .Y(new_n1476_));
  NAND2X1  g0995(.A(new_n1476_), .B(\V1481(0) ), .Y(new_n1477_));
  NOR3X1   g0996(.A(\V149(2) ), .B(new_n483_), .C(new_n497_), .Y(new_n1478_));
  OR4X1    g0997(.A(new_n1047_), .B(new_n498_), .C(\V149(4) ), .D(\V149(6) ), .Y(new_n1479_));
  NAND3X1  g0998(.A(new_n485_), .B(\V149(4) ), .C(new_n501_), .Y(new_n1480_));
  OR4X1    g0999(.A(new_n1480_), .B(new_n498_), .C(new_n527_), .D(\V149(6) ), .Y(new_n1481_));
  NOR4X1   g1000(.A(new_n718_), .B(new_n498_), .C(\V149(4) ), .D(new_n495_), .Y(new_n1482_));
  INVX1    g1001(.A(new_n1482_), .Y(new_n1483_));
  NAND3X1  g1002(.A(\V149(3) ), .B(new_n527_), .C(\V149(7) ), .Y(new_n1484_));
  NOR4X1   g1003(.A(new_n1484_), .B(new_n498_), .C(\V149(4) ), .D(\V149(6) ), .Y(new_n1485_));
  NOR4X1   g1004(.A(new_n1485_), .B(new_n719_), .C(new_n498_), .D(new_n485_), .Y(new_n1486_));
  NAND2X1  g1005(.A(new_n1486_), .B(new_n1483_), .Y(new_n1487_));
  NAND3X1  g1006(.A(new_n1487_), .B(new_n1481_), .C(new_n1479_), .Y(new_n1488_));
  NOR3X1   g1007(.A(new_n484_), .B(new_n483_), .C(new_n497_), .Y(new_n1489_));
  NOR3X1   g1008(.A(new_n484_), .B(\V149(1) ), .C(new_n497_), .Y(new_n1490_));
  NOR4X1   g1009(.A(new_n1490_), .B(new_n1489_), .C(new_n1488_), .D(new_n1478_), .Y(new_n1491_));
  AND2X1   g1010(.A(new_n1488_), .B(\V1864(0) ), .Y(new_n1492_));
  NOR3X1   g1011(.A(new_n1492_), .B(new_n1491_), .C(new_n578_), .Y(new_n1493_));
  OR2X1    g1012(.A(new_n1493_), .B(new_n1096_), .Y(new_n1494_));
  OR4X1    g1013(.A(new_n1494_), .B(new_n1477_), .C(new_n1473_), .D(new_n1431_), .Y(\V798(0) ));
  AND2X1   g1014(.A(new_n504_), .B(new_n492_), .Y(V801));
  INVX1    g1015(.A(\V279(0) ), .Y(new_n1497_));
  NOR2X1   g1016(.A(new_n559_), .B(new_n493_), .Y(new_n1498_));
  MX2X1    g1017(.A(new_n1497_), .B(\V149(5) ), .S0(new_n1498_), .Y(\V821(0) ));
  OAI21X1  g1018(.A0(new_n559_), .A1(new_n493_), .B0(new_n1497_), .Y(new_n1500_));
  INVX1    g1019(.A(\V280(0) ), .Y(new_n1501_));
  NOR3X1   g1020(.A(new_n1498_), .B(new_n1501_), .C(new_n1497_), .Y(new_n1502_));
  AOI21X1  g1021(.A0(new_n1498_), .A1(\V149(4) ), .B0(new_n1502_), .Y(new_n1503_));
  OAI21X1  g1022(.A0(new_n1500_), .A1(\V280(0) ), .B0(new_n1503_), .Y(\V826(0) ));
  NOR2X1   g1023(.A(new_n1493_), .B(new_n493_), .Y(new_n1505_));
  AND2X1   g1024(.A(new_n1488_), .B(\V56(0) ), .Y(new_n1506_));
  INVX1    g1025(.A(new_n492_), .Y(new_n1507_));
  NOR2X1   g1026(.A(new_n504_), .B(new_n1507_), .Y(new_n1508_));
  NOR4X1   g1027(.A(new_n1441_), .B(new_n572_), .C(new_n504_), .D(new_n531_), .Y(new_n1509_));
  NOR4X1   g1028(.A(new_n1509_), .B(new_n1508_), .C(new_n1506_), .D(new_n1505_), .Y(new_n1510_));
  NOR3X1   g1029(.A(new_n1510_), .B(new_n1475_), .C(new_n1096_), .Y(V966));
  INVX1    g1030(.A(new_n1104_), .Y(new_n1512_));
  NOR4X1   g1031(.A(new_n562_), .B(new_n1102_), .C(new_n524_), .D(new_n486_), .Y(new_n1513_));
  AOI21X1  g1032(.A0(new_n1513_), .A1(new_n1512_), .B0(new_n1005_), .Y(new_n1514_));
  AOI21X1  g1033(.A0(new_n577_), .A1(new_n576_), .B0(new_n1001_), .Y(new_n1515_));
  INVX1    g1034(.A(new_n1467_), .Y(new_n1516_));
  NOR4X1   g1035(.A(new_n1509_), .B(new_n1488_), .C(new_n1516_), .D(new_n531_), .Y(new_n1517_));
  NOR3X1   g1036(.A(new_n1517_), .B(new_n1515_), .C(new_n1514_), .Y(new_n1518_));
  NOR3X1   g1037(.A(new_n1518_), .B(new_n1475_), .C(new_n1096_), .Y(V986));
  INVX1    g1038(.A(new_n1315_), .Y(\V1243(3) ));
  INVX1    g1039(.A(new_n1335_), .Y(\V1243(2) ));
  INVX1    g1040(.A(new_n1355_), .Y(\V1243(1) ));
  INVX1    g1041(.A(\V2(0) ), .Y(new_n1523_));
  NOR3X1   g1042(.A(new_n1523_), .B(\V13(0) ), .C(new_n1435_), .Y(V1256));
  OR2X1    g1043(.A(\V63(0) ), .B(\V60(0) ), .Y(new_n1525_));
  AND2X1   g1044(.A(new_n1525_), .B(new_n529_), .Y(new_n1526_));
  NOR3X1   g1045(.A(new_n1006_), .B(new_n562_), .C(new_n557_), .Y(new_n1527_));
  AND2X1   g1046(.A(new_n994_), .B(new_n559_), .Y(new_n1528_));
  AND2X1   g1047(.A(new_n1528_), .B(new_n554_), .Y(new_n1529_));
  AOI21X1  g1048(.A0(new_n1529_), .A1(new_n1527_), .B0(new_n532_), .Y(new_n1530_));
  AND2X1   g1049(.A(new_n1049_), .B(new_n532_), .Y(new_n1531_));
  OR4X1    g1050(.A(new_n1531_), .B(new_n1523_), .C(new_n1438_), .D(\V174(0) ), .Y(new_n1532_));
  NOR4X1   g1051(.A(new_n1532_), .B(new_n1530_), .C(new_n1526_), .D(\V35(0) ), .Y(V1257));
  AND2X1   g1052(.A(\V3(0) ), .B(\V9(0) ), .Y(V1259));
  AND2X1   g1053(.A(\V3(0) ), .B(\V11(0) ), .Y(V1260));
  AND2X1   g1054(.A(V1260), .B(new_n1001_), .Y(V1261));
  NOR3X1   g1055(.A(new_n1448_), .B(\V13(0) ), .C(new_n1435_), .Y(V1262));
  AND2X1   g1056(.A(\V4(0) ), .B(\V9(0) ), .Y(V1263));
  AND2X1   g1057(.A(\V4(0) ), .B(\V12(0) ), .Y(V1264));
  AND2X1   g1058(.A(V1264), .B(\V52(0) ), .Y(V1265));
  AND2X1   g1059(.A(\V4(0) ), .B(\V11(0) ), .Y(V1266));
  AND2X1   g1060(.A(\V2(0) ), .B(\V11(0) ), .Y(V1267));
  NAND4X1  g1061(.A(new_n1432_), .B(new_n537_), .C(\V14(0) ), .D(\V62(0) ), .Y(new_n1543_));
  NOR2X1   g1062(.A(new_n503_), .B(\V174(0) ), .Y(new_n1544_));
  OR4X1    g1063(.A(new_n1104_), .B(new_n993_), .C(new_n562_), .D(new_n486_), .Y(new_n1545_));
  OR4X1    g1064(.A(new_n1545_), .B(new_n995_), .C(new_n1102_), .D(new_n524_), .Y(new_n1546_));
  NAND3X1  g1065(.A(new_n1415_), .B(new_n922_), .C(\V59(0) ), .Y(new_n1547_));
  NOR4X1   g1066(.A(new_n1547_), .B(new_n1546_), .C(new_n1544_), .D(new_n719_), .Y(new_n1548_));
  NAND3X1  g1067(.A(new_n1548_), .B(new_n1432_), .C(\V14(0) ), .Y(new_n1549_));
  NAND2X1  g1068(.A(new_n1549_), .B(new_n1543_), .Y(\V1274(0) ));
  INVX1    g1069(.A(new_n507_), .Y(new_n1551_));
  NOR3X1   g1070(.A(new_n536_), .B(new_n535_), .C(new_n534_), .Y(new_n1552_));
  OAI22X1  g1071(.A0(new_n564_), .A1(\V302(0) ), .B0(new_n500_), .B1(\V174(0) ), .Y(new_n1553_));
  NOR3X1   g1072(.A(new_n1553_), .B(new_n1552_), .C(new_n1420_), .Y(new_n1554_));
  OR2X1    g1073(.A(new_n1096_), .B(\V289(0) ), .Y(new_n1555_));
  NOR4X1   g1074(.A(new_n1555_), .B(new_n1554_), .C(new_n1029_), .D(new_n920_), .Y(new_n1556_));
  NOR4X1   g1075(.A(new_n1556_), .B(new_n1029_), .C(new_n920_), .D(new_n1551_), .Y(new_n1557_));
  AND2X1   g1076(.A(new_n1453_), .B(new_n507_), .Y(new_n1558_));
  AOI21X1  g1077(.A0(new_n1557_), .A1(new_n503_), .B0(new_n1558_), .Y(new_n1559_));
  AOI21X1  g1078(.A0(new_n1458_), .A1(\V56(0) ), .B0(new_n1096_), .Y(new_n1560_));
  AND2X1   g1079(.A(new_n1560_), .B(\V213(0) ), .Y(new_n1561_));
  OR4X1    g1080(.A(\V165(3) ), .B(\V165(7) ), .C(\V165(5) ), .D(\V165(4) ), .Y(new_n1562_));
  OAI22X1  g1081(.A0(new_n1562_), .A1(\V165(6) ), .B0(new_n1027_), .B1(new_n1026_), .Y(new_n1563_));
  MX2X1    g1082(.A(new_n1563_), .B(new_n1561_), .S0(new_n1559_), .Y(\V1281(0) ));
  AND2X1   g1083(.A(new_n1560_), .B(\V213(5) ), .Y(new_n1565_));
  MX2X1    g1084(.A(new_n1565_), .B(\V165(7) ), .S0(new_n1558_), .Y(\V1297(4) ));
  AND2X1   g1085(.A(new_n1560_), .B(\V213(4) ), .Y(new_n1567_));
  MX2X1    g1086(.A(new_n1567_), .B(\V165(6) ), .S0(new_n1558_), .Y(\V1297(3) ));
  AND2X1   g1087(.A(new_n1560_), .B(\V213(3) ), .Y(new_n1569_));
  MX2X1    g1088(.A(new_n1569_), .B(\V165(5) ), .S0(new_n1558_), .Y(\V1297(2) ));
  AND2X1   g1089(.A(new_n1560_), .B(\V213(2) ), .Y(new_n1571_));
  MX2X1    g1090(.A(new_n1571_), .B(\V165(4) ), .S0(new_n1558_), .Y(\V1297(1) ));
  AND2X1   g1091(.A(new_n1560_), .B(\V213(1) ), .Y(new_n1573_));
  MX2X1    g1092(.A(new_n1573_), .B(\V165(3) ), .S0(new_n1558_), .Y(\V1297(0) ));
  OR4X1    g1093(.A(new_n1475_), .B(new_n1420_), .C(new_n1049_), .D(new_n1096_), .Y(new_n1575_));
  OR4X1    g1094(.A(new_n1575_), .B(new_n1008_), .C(new_n1007_), .D(new_n578_), .Y(new_n1576_));
  NOR4X1   g1095(.A(new_n1576_), .B(new_n1069_), .C(new_n1006_), .D(new_n1001_), .Y(V1365));
  INVX1    g1096(.A(\V268(5) ), .Y(V1375));
  INVX1    g1097(.A(V782), .Y(new_n1579_));
  NOR3X1   g1098(.A(new_n1579_), .B(new_n1410_), .C(new_n493_), .Y(V1378));
  NOR4X1   g1099(.A(new_n1405_), .B(new_n580_), .C(\V802(0) ), .D(\V248(0) ), .Y(new_n1581_));
  NAND3X1  g1100(.A(new_n1581_), .B(new_n1234_), .C(new_n524_), .Y(new_n1582_));
  NAND2X1  g1101(.A(new_n493_), .B(\V248(0) ), .Y(new_n1583_));
  AND2X1   g1102(.A(new_n580_), .B(new_n493_), .Y(new_n1584_));
  NOR2X1   g1103(.A(new_n1234_), .B(\V802(0) ), .Y(new_n1585_));
  NOR4X1   g1104(.A(new_n1585_), .B(new_n1584_), .C(new_n1405_), .D(new_n1410_), .Y(new_n1586_));
  AOI21X1  g1105(.A0(new_n1586_), .A1(new_n1583_), .B0(new_n1238_), .Y(new_n1587_));
  AOI21X1  g1106(.A0(new_n1587_), .A1(new_n1582_), .B0(new_n1579_), .Y(V1380));
  OR2X1    g1107(.A(\V13(0) ), .B(new_n1435_), .Y(new_n1589_));
  AOI21X1  g1108(.A0(new_n536_), .A1(new_n564_), .B0(new_n493_), .Y(new_n1590_));
  OAI21X1  g1109(.A0(new_n1590_), .A1(new_n1102_), .B0(\V7(0) ), .Y(new_n1591_));
  NOR2X1   g1110(.A(new_n1591_), .B(new_n1589_), .Y(V1382));
  NAND4X1  g1111(.A(new_n1055_), .B(new_n1048_), .C(new_n1018_), .D(\V56(0) ), .Y(new_n1593_));
  NOR3X1   g1112(.A(new_n1593_), .B(new_n1589_), .C(new_n1443_), .Y(V1384));
  NOR3X1   g1113(.A(\V50(0) ), .B(\V62(0) ), .C(\V56(0) ), .Y(new_n1595_));
  NOR4X1   g1114(.A(new_n1595_), .B(new_n1589_), .C(new_n595_), .D(new_n1443_), .Y(V1386));
  OR4X1    g1115(.A(new_n1475_), .B(new_n572_), .C(new_n1096_), .D(\V165(5) ), .Y(new_n1597_));
  OR4X1    g1116(.A(new_n1597_), .B(new_n490_), .C(new_n488_), .D(\V165(4) ), .Y(new_n1598_));
  NAND4X1  g1117(.A(new_n1432_), .B(new_n1098_), .C(\V14(0) ), .D(\V65(0) ), .Y(new_n1599_));
  OAI22X1  g1118(.A0(new_n1599_), .A1(new_n555_), .B0(new_n1598_), .B1(new_n489_), .Y(\V1392(0) ));
  INVX1    g1119(.A(\V1(0) ), .Y(new_n1601_));
  NOR3X1   g1120(.A(new_n1601_), .B(\V13(0) ), .C(new_n1435_), .Y(V1426));
  AND2X1   g1121(.A(\V11(0) ), .B(\V1(0) ), .Y(V1428));
  AND2X1   g1122(.A(\V12(0) ), .B(\V1(0) ), .Y(V1429));
  NOR3X1   g1123(.A(new_n905_), .B(new_n1447_), .C(new_n1601_), .Y(V1431));
  NOR3X1   g1124(.A(new_n1475_), .B(new_n1096_), .C(new_n991_), .Y(V1432));
  INVX1    g1125(.A(\V277(0) ), .Y(new_n1607_));
  NOR3X1   g1126(.A(new_n562_), .B(new_n1607_), .C(new_n1096_), .Y(new_n1608_));
  OR2X1    g1127(.A(new_n1608_), .B(new_n1464_), .Y(\V1439(0) ));
  OR2X1    g1128(.A(new_n580_), .B(new_n1096_), .Y(\V1440(0) ));
  INVX1    g1129(.A(\V268(0) ), .Y(new_n1611_));
  INVX1    g1130(.A(\V268(1) ), .Y(new_n1612_));
  INVX1    g1131(.A(\V268(2) ), .Y(new_n1613_));
  INVX1    g1132(.A(\V268(4) ), .Y(new_n1614_));
  NAND2X1  g1133(.A(\V268(3) ), .B(\V268(5) ), .Y(new_n1615_));
  NOR4X1   g1134(.A(new_n1615_), .B(new_n1614_), .C(new_n1613_), .D(new_n1612_), .Y(new_n1616_));
  INVX1    g1135(.A(new_n1616_), .Y(new_n1617_));
  OAI22X1  g1136(.A0(new_n1617_), .A1(new_n1611_), .B0(new_n1595_), .B1(new_n595_), .Y(new_n1618_));
  NOR2X1   g1137(.A(new_n1618_), .B(new_n1096_), .Y(new_n1619_));
  AND2X1   g1138(.A(new_n1618_), .B(\V14(0) ), .Y(new_n1620_));
  MX2X1    g1139(.A(new_n1620_), .B(new_n1619_), .S0(\V258(0) ), .Y(\V1451(0) ));
  INVX1    g1140(.A(\V259(0) ), .Y(new_n1622_));
  NOR3X1   g1141(.A(new_n1595_), .B(new_n595_), .C(\V258(0) ), .Y(new_n1623_));
  NOR3X1   g1142(.A(new_n1617_), .B(new_n1611_), .C(new_n1461_), .Y(new_n1624_));
  OR4X1    g1143(.A(new_n1624_), .B(new_n1623_), .C(new_n1622_), .D(new_n1096_), .Y(new_n1625_));
  OAI21X1  g1144(.A0(new_n1624_), .A1(new_n1623_), .B0(new_n1622_), .Y(new_n1626_));
  OAI21X1  g1145(.A0(new_n1626_), .A1(new_n1096_), .B0(new_n1625_), .Y(\V1459(0) ));
  NOR4X1   g1146(.A(new_n1595_), .B(new_n595_), .C(\V259(0) ), .D(\V258(0) ), .Y(new_n1628_));
  AOI21X1  g1147(.A0(new_n1624_), .A1(\V259(0) ), .B0(new_n1628_), .Y(new_n1629_));
  NAND3X1  g1148(.A(new_n1629_), .B(\V260(0) ), .C(\V14(0) ), .Y(new_n1630_));
  OR2X1    g1149(.A(new_n1629_), .B(\V260(0) ), .Y(new_n1631_));
  OAI21X1  g1150(.A0(new_n1631_), .A1(new_n1096_), .B0(new_n1630_), .Y(\V1467(0) ));
  NOR4X1   g1151(.A(new_n1475_), .B(new_n1075_), .C(new_n1417_), .D(new_n1096_), .Y(V1470));
  OAI21X1  g1152(.A0(new_n1021_), .A1(new_n1020_), .B0(new_n564_), .Y(new_n1634_));
  NAND3X1  g1153(.A(\V1757(0) ), .B(new_n1051_), .C(\V802(0) ), .Y(new_n1635_));
  NAND3X1  g1154(.A(new_n1635_), .B(new_n1634_), .C(new_n1055_), .Y(\V1480(0) ));
  INVX1    g1155(.A(\V216(0) ), .Y(new_n1637_));
  OR4X1    g1156(.A(\V69(0) ), .B(\V68(0) ), .C(\V70(0) ), .D(\V66(0) ), .Y(new_n1638_));
  NAND4X1  g1157(.A(new_n1638_), .B(new_n1426_), .C(\V14(0) ), .D(\V215(0) ), .Y(new_n1639_));
  OAI21X1  g1158(.A0(new_n1637_), .A1(\V214(0) ), .B0(new_n1639_), .Y(\V1492(0) ));
  INVX1    g1159(.A(\V175(0) ), .Y(\V1495(0) ));
  NOR4X1   g1160(.A(new_n484_), .B(\V149(1) ), .C(\V149(0) ), .D(new_n531_), .Y(new_n1642_));
  AOI22X1  g1161(.A0(new_n1642_), .A1(\V149(7) ), .B0(new_n1028_), .B1(new_n1051_), .Y(new_n1643_));
  NAND3X1  g1162(.A(new_n996_), .B(new_n1418_), .C(\V56(0) ), .Y(new_n1644_));
  NOR2X1   g1163(.A(\V274(0) ), .B(\V271(0) ), .Y(new_n1645_));
  INVX1    g1164(.A(\V177(0) ), .Y(new_n1646_));
  INVX1    g1165(.A(\V171(0) ), .Y(new_n1647_));
  OR2X1    g1166(.A(new_n535_), .B(new_n531_), .Y(new_n1648_));
  OAI22X1  g1167(.A0(new_n1648_), .A1(new_n1647_), .B0(new_n589_), .B1(new_n561_), .Y(new_n1649_));
  NOR4X1   g1168(.A(new_n1649_), .B(new_n1027_), .C(new_n1646_), .D(\V248(0) ), .Y(new_n1650_));
  NOR3X1   g1169(.A(new_n1650_), .B(new_n1645_), .C(new_n1116_), .Y(new_n1651_));
  NAND2X1  g1170(.A(new_n1651_), .B(new_n1644_), .Y(new_n1652_));
  NAND3X1  g1171(.A(new_n1652_), .B(new_n1643_), .C(new_n1428_), .Y(\V1536(0) ));
  OR4X1    g1172(.A(new_n868_), .B(new_n866_), .C(new_n860_), .D(new_n854_), .Y(new_n1654_));
  OR4X1    g1173(.A(new_n1654_), .B(new_n767_), .C(new_n759_), .D(new_n748_), .Y(new_n1655_));
  OR2X1    g1174(.A(new_n1655_), .B(new_n732_), .Y(new_n1656_));
  MX2X1    g1175(.A(new_n1656_), .B(new_n1428_), .S0(\V1536(0) ), .Y(\V1512(3) ));
  INVX1    g1176(.A(new_n1440_), .Y(new_n1658_));
  INVX1    g1177(.A(new_n1643_), .Y(new_n1659_));
  NAND3X1  g1178(.A(new_n1659_), .B(new_n1658_), .C(new_n1428_), .Y(new_n1660_));
  OR2X1    g1179(.A(new_n896_), .B(new_n854_), .Y(new_n1661_));
  OR4X1    g1180(.A(new_n1661_), .B(new_n883_), .C(new_n866_), .D(new_n789_), .Y(new_n1662_));
  OR4X1    g1181(.A(new_n1662_), .B(new_n845_), .C(new_n759_), .D(new_n732_), .Y(new_n1663_));
  MX2X1    g1182(.A(new_n1663_), .B(new_n1660_), .S0(\V1536(0) ), .Y(\V1512(2) ));
  NAND2X1  g1183(.A(new_n1440_), .B(new_n1428_), .Y(new_n1665_));
  OR4X1    g1184(.A(new_n1661_), .B(new_n890_), .C(new_n860_), .D(new_n816_), .Y(new_n1666_));
  OR4X1    g1185(.A(new_n1666_), .B(new_n845_), .C(new_n748_), .D(new_n732_), .Y(new_n1667_));
  MX2X1    g1186(.A(new_n1667_), .B(new_n1665_), .S0(\V1536(0) ), .Y(\V1512(1) ));
  AND2X1   g1187(.A(new_n1432_), .B(\V68(0) ), .Y(new_n1669_));
  AND2X1   g1188(.A(new_n1669_), .B(\V14(0) ), .Y(V1537));
  OAI21X1  g1189(.A0(\V50(0) ), .A1(\V69(0) ), .B0(new_n1432_), .Y(new_n1671_));
  NOR2X1   g1190(.A(new_n1671_), .B(new_n1096_), .Y(V1539));
  INVX1    g1191(.A(new_n1590_), .Y(new_n1673_));
  OR4X1    g1192(.A(new_n564_), .B(\V802(0) ), .C(\V239(4) ), .D(new_n485_), .Y(new_n1674_));
  OAI21X1  g1193(.A0(new_n559_), .A1(\V802(0) ), .B0(\V1243(9) ), .Y(new_n1675_));
  OAI21X1  g1194(.A0(new_n1675_), .A1(new_n1673_), .B0(new_n1674_), .Y(\V1552(1) ));
  XOR2X1   g1195(.A(\V239(3) ), .B(new_n933_), .Y(new_n1677_));
  OR4X1    g1196(.A(new_n1677_), .B(new_n1590_), .C(new_n559_), .D(\V802(0) ), .Y(new_n1678_));
  OAI21X1  g1197(.A0(new_n559_), .A1(\V802(0) ), .B0(\V1243(8) ), .Y(new_n1679_));
  OAI21X1  g1198(.A0(new_n1679_), .A1(new_n1673_), .B0(new_n1678_), .Y(\V1552(0) ));
  INVX1    g1199(.A(new_n1459_), .Y(new_n1681_));
  NAND4X1  g1200(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(1) ), .Y(new_n1682_));
  AND2X1   g1201(.A(new_n1463_), .B(\V132(0) ), .Y(new_n1683_));
  AND2X1   g1202(.A(new_n1683_), .B(new_n1681_), .Y(new_n1684_));
  INVX1    g1203(.A(\V108(5) ), .Y(new_n1685_));
  NOR3X1   g1204(.A(new_n1463_), .B(new_n1459_), .C(new_n1685_), .Y(new_n1686_));
  MX2X1    g1205(.A(new_n1684_), .B(new_n1686_), .S0(new_n1482_), .Y(\V1953(0) ));
  XOR2X1   g1206(.A(\V1953(0) ), .B(new_n1682_), .Y(new_n1688_));
  INVX1    g1207(.A(new_n1458_), .Y(new_n1689_));
  INVX1    g1208(.A(new_n1460_), .Y(new_n1690_));
  NAND4X1  g1209(.A(new_n1463_), .B(new_n1690_), .C(new_n1689_), .D(\V124(5) ), .Y(new_n1691_));
  NOR2X1   g1210(.A(new_n1691_), .B(new_n1485_), .Y(new_n1692_));
  INVX1    g1211(.A(new_n1463_), .Y(new_n1693_));
  NAND4X1  g1212(.A(new_n1693_), .B(new_n1460_), .C(new_n1689_), .D(\V100(5) ), .Y(new_n1694_));
  INVX1    g1213(.A(\V213(5) ), .Y(new_n1695_));
  OR4X1    g1214(.A(new_n1463_), .B(new_n1460_), .C(new_n1689_), .D(new_n1695_), .Y(new_n1696_));
  AOI21X1  g1215(.A0(new_n1696_), .A1(new_n1694_), .B0(new_n1485_), .Y(new_n1697_));
  OR2X1    g1216(.A(new_n1697_), .B(new_n1692_), .Y(\V1921(5) ));
  INVX1    g1217(.A(new_n1485_), .Y(new_n1699_));
  INVX1    g1218(.A(\V124(4) ), .Y(new_n1700_));
  NOR4X1   g1219(.A(new_n1693_), .B(new_n1460_), .C(new_n1458_), .D(new_n1700_), .Y(new_n1701_));
  INVX1    g1220(.A(\V108(4) ), .Y(new_n1702_));
  NOR4X1   g1221(.A(new_n1463_), .B(new_n1460_), .C(new_n1458_), .D(new_n1702_), .Y(new_n1703_));
  MX2X1    g1222(.A(new_n1703_), .B(new_n1701_), .S0(new_n1699_), .Y(new_n1704_));
  NAND4X1  g1223(.A(new_n1693_), .B(new_n1460_), .C(new_n1689_), .D(\V100(4) ), .Y(new_n1705_));
  NAND4X1  g1224(.A(new_n1693_), .B(new_n1690_), .C(new_n1458_), .D(\V213(4) ), .Y(new_n1706_));
  AOI21X1  g1225(.A0(new_n1706_), .A1(new_n1705_), .B0(new_n1485_), .Y(new_n1707_));
  NOR2X1   g1226(.A(new_n1707_), .B(new_n1704_), .Y(new_n1708_));
  XOR2X1   g1227(.A(new_n1708_), .B(\V1921(5) ), .Y(new_n1709_));
  XOR2X1   g1228(.A(new_n1709_), .B(new_n1688_), .Y(new_n1710_));
  INVX1    g1229(.A(\V124(3) ), .Y(new_n1711_));
  NOR4X1   g1230(.A(new_n1693_), .B(new_n1460_), .C(new_n1458_), .D(new_n1711_), .Y(new_n1712_));
  INVX1    g1231(.A(\V108(3) ), .Y(new_n1713_));
  NOR4X1   g1232(.A(new_n1463_), .B(new_n1460_), .C(new_n1458_), .D(new_n1713_), .Y(new_n1714_));
  MX2X1    g1233(.A(new_n1714_), .B(new_n1712_), .S0(new_n1699_), .Y(new_n1715_));
  NAND4X1  g1234(.A(new_n1693_), .B(new_n1460_), .C(new_n1689_), .D(\V100(3) ), .Y(new_n1716_));
  NAND4X1  g1235(.A(new_n1693_), .B(new_n1690_), .C(new_n1458_), .D(\V213(3) ), .Y(new_n1717_));
  AOI21X1  g1236(.A0(new_n1717_), .A1(new_n1716_), .B0(new_n1485_), .Y(new_n1718_));
  NOR2X1   g1237(.A(new_n1718_), .B(new_n1715_), .Y(new_n1719_));
  INVX1    g1238(.A(\V124(2) ), .Y(new_n1720_));
  NOR4X1   g1239(.A(new_n1693_), .B(new_n1460_), .C(new_n1458_), .D(new_n1720_), .Y(new_n1721_));
  INVX1    g1240(.A(\V108(2) ), .Y(new_n1722_));
  NOR4X1   g1241(.A(new_n1463_), .B(new_n1460_), .C(new_n1458_), .D(new_n1722_), .Y(new_n1723_));
  MX2X1    g1242(.A(new_n1723_), .B(new_n1721_), .S0(new_n1699_), .Y(new_n1724_));
  NAND4X1  g1243(.A(new_n1693_), .B(new_n1460_), .C(new_n1689_), .D(\V100(2) ), .Y(new_n1725_));
  NAND4X1  g1244(.A(new_n1693_), .B(new_n1690_), .C(new_n1458_), .D(\V213(2) ), .Y(new_n1726_));
  AOI21X1  g1245(.A0(new_n1726_), .A1(new_n1725_), .B0(new_n1485_), .Y(new_n1727_));
  NOR2X1   g1246(.A(new_n1727_), .B(new_n1724_), .Y(new_n1728_));
  XOR2X1   g1247(.A(new_n1728_), .B(new_n1719_), .Y(new_n1729_));
  INVX1    g1248(.A(\V124(1) ), .Y(new_n1730_));
  NOR4X1   g1249(.A(new_n1693_), .B(new_n1460_), .C(new_n1458_), .D(new_n1730_), .Y(new_n1731_));
  INVX1    g1250(.A(\V108(1) ), .Y(new_n1732_));
  NOR4X1   g1251(.A(new_n1463_), .B(new_n1460_), .C(new_n1458_), .D(new_n1732_), .Y(new_n1733_));
  MX2X1    g1252(.A(new_n1733_), .B(new_n1731_), .S0(new_n1699_), .Y(new_n1734_));
  NAND4X1  g1253(.A(new_n1693_), .B(new_n1460_), .C(new_n1689_), .D(\V100(1) ), .Y(new_n1735_));
  NAND4X1  g1254(.A(new_n1693_), .B(new_n1690_), .C(new_n1458_), .D(\V213(1) ), .Y(new_n1736_));
  AOI21X1  g1255(.A0(new_n1736_), .A1(new_n1735_), .B0(new_n1485_), .Y(new_n1737_));
  OR2X1    g1256(.A(new_n1737_), .B(new_n1734_), .Y(\V1921(1) ));
  INVX1    g1257(.A(\V124(0) ), .Y(new_n1739_));
  NOR4X1   g1258(.A(new_n1693_), .B(new_n1460_), .C(new_n1458_), .D(new_n1739_), .Y(new_n1740_));
  INVX1    g1259(.A(\V108(0) ), .Y(new_n1741_));
  NOR4X1   g1260(.A(new_n1463_), .B(new_n1460_), .C(new_n1458_), .D(new_n1741_), .Y(new_n1742_));
  MX2X1    g1261(.A(new_n1742_), .B(new_n1740_), .S0(new_n1699_), .Y(new_n1743_));
  NAND4X1  g1262(.A(new_n1693_), .B(new_n1460_), .C(new_n1689_), .D(\V100(0) ), .Y(new_n1744_));
  NAND4X1  g1263(.A(new_n1693_), .B(new_n1690_), .C(new_n1458_), .D(\V213(0) ), .Y(new_n1745_));
  AOI21X1  g1264(.A0(new_n1745_), .A1(new_n1744_), .B0(new_n1485_), .Y(new_n1746_));
  NOR2X1   g1265(.A(new_n1746_), .B(new_n1743_), .Y(new_n1747_));
  XOR2X1   g1266(.A(new_n1747_), .B(\V1921(1) ), .Y(new_n1748_));
  XOR2X1   g1267(.A(new_n1748_), .B(new_n1729_), .Y(new_n1749_));
  XOR2X1   g1268(.A(new_n1749_), .B(new_n1710_), .Y(\V1613(0) ));
  AND2X1   g1269(.A(new_n1459_), .B(\V118(7) ), .Y(new_n1751_));
  AND2X1   g1270(.A(new_n1681_), .B(\V46(0) ), .Y(new_n1752_));
  MX2X1    g1271(.A(new_n1752_), .B(new_n1751_), .S0(new_n1099_), .Y(\V1960(1) ));
  AND2X1   g1272(.A(new_n1459_), .B(\V118(6) ), .Y(new_n1754_));
  AND2X1   g1273(.A(new_n1681_), .B(\V48(0) ), .Y(new_n1755_));
  MX2X1    g1274(.A(new_n1755_), .B(new_n1754_), .S0(new_n1099_), .Y(\V1960(0) ));
  XOR2X1   g1275(.A(\V1960(0) ), .B(\V1960(1) ), .Y(new_n1757_));
  NAND4X1  g1276(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(7) ), .Y(new_n1758_));
  NAND4X1  g1277(.A(new_n1483_), .B(new_n1693_), .C(new_n1459_), .D(\V118(5) ), .Y(new_n1759_));
  NAND2X1  g1278(.A(new_n1759_), .B(new_n1758_), .Y(\V1953(7) ));
  NAND4X1  g1279(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(6) ), .Y(new_n1761_));
  NAND4X1  g1280(.A(new_n1483_), .B(new_n1693_), .C(new_n1459_), .D(\V118(4) ), .Y(new_n1762_));
  NAND2X1  g1281(.A(new_n1762_), .B(new_n1761_), .Y(\V1953(6) ));
  XOR2X1   g1282(.A(\V1953(6) ), .B(\V1953(7) ), .Y(new_n1764_));
  XOR2X1   g1283(.A(new_n1764_), .B(new_n1757_), .Y(new_n1765_));
  NAND4X1  g1284(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(5) ), .Y(new_n1766_));
  NAND4X1  g1285(.A(new_n1483_), .B(new_n1693_), .C(new_n1459_), .D(\V118(3) ), .Y(new_n1767_));
  NAND2X1  g1286(.A(new_n1767_), .B(new_n1766_), .Y(\V1953(5) ));
  NAND4X1  g1287(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(4) ), .Y(new_n1769_));
  NAND4X1  g1288(.A(new_n1483_), .B(new_n1693_), .C(new_n1459_), .D(\V118(2) ), .Y(new_n1770_));
  NAND2X1  g1289(.A(new_n1770_), .B(new_n1769_), .Y(\V1953(4) ));
  XOR2X1   g1290(.A(\V1953(4) ), .B(\V1953(5) ), .Y(new_n1772_));
  NAND4X1  g1291(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(3) ), .Y(new_n1773_));
  NAND4X1  g1292(.A(new_n1483_), .B(new_n1693_), .C(new_n1459_), .D(\V118(1) ), .Y(new_n1774_));
  AND2X1   g1293(.A(new_n1774_), .B(new_n1773_), .Y(new_n1775_));
  NAND4X1  g1294(.A(new_n1483_), .B(new_n1463_), .C(new_n1681_), .D(\V132(2) ), .Y(new_n1776_));
  NAND4X1  g1295(.A(new_n1483_), .B(new_n1693_), .C(new_n1459_), .D(\V118(0) ), .Y(new_n1777_));
  NAND2X1  g1296(.A(new_n1777_), .B(new_n1776_), .Y(\V1953(2) ));
  XOR2X1   g1297(.A(\V1953(2) ), .B(new_n1775_), .Y(new_n1779_));
  XOR2X1   g1298(.A(new_n1779_), .B(new_n1772_), .Y(new_n1780_));
  XOR2X1   g1299(.A(new_n1780_), .B(new_n1765_), .Y(\V1613(1) ));
  AOI22X1  g1300(.A0(new_n1429_), .A1(\V174(0) ), .B0(\V292(0) ), .B1(\V1864(0) ), .Y(new_n1782_));
  AOI22X1  g1301(.A0(new_n920_), .A1(\V174(0) ), .B0(new_n491_), .B1(new_n488_), .Y(new_n1783_));
  NAND2X1  g1302(.A(new_n1783_), .B(new_n1782_), .Y(\V1620(0) ));
  OR2X1    g1303(.A(new_n1067_), .B(\V294(0) ), .Y(new_n1785_));
  AND2X1   g1304(.A(\V91(1) ), .B(\V62(0) ), .Y(new_n1786_));
  AND2X1   g1305(.A(\V91(0) ), .B(\V59(0) ), .Y(new_n1787_));
  OR2X1    g1306(.A(new_n1787_), .B(new_n1786_), .Y(new_n1788_));
  AOI21X1  g1307(.A0(new_n1788_), .A1(new_n1049_), .B0(new_n1396_), .Y(new_n1789_));
  OAI21X1  g1308(.A0(new_n1785_), .A1(new_n1105_), .B0(new_n1789_), .Y(\V1629(0) ));
  NOR2X1   g1309(.A(new_n1066_), .B(new_n501_), .Y(new_n1791_));
  OR2X1    g1310(.A(new_n1791_), .B(new_n1556_), .Y(new_n1792_));
  OR2X1    g1311(.A(new_n1792_), .B(new_n1078_), .Y(\V1645(0) ));
  NOR2X1   g1312(.A(new_n1086_), .B(new_n583_), .Y(new_n1794_));
  NOR4X1   g1313(.A(new_n1794_), .B(new_n578_), .C(\V249(0) ), .D(\V289(0) ), .Y(new_n1795_));
  NAND3X1  g1314(.A(new_n1795_), .B(\V295(0) ), .C(new_n1452_), .Y(\V1652(0) ));
  INVX1    g1315(.A(\V289(0) ), .Y(new_n1797_));
  NAND2X1  g1316(.A(new_n988_), .B(new_n1797_), .Y(new_n1798_));
  NOR2X1   g1317(.A(new_n1798_), .B(\V802(0) ), .Y(new_n1799_));
  NOR4X1   g1318(.A(\V260(0) ), .B(\V259(0) ), .C(new_n1461_), .D(\V59(0) ), .Y(new_n1800_));
  NAND2X1  g1319(.A(\V262(0) ), .B(\V14(0) ), .Y(new_n1801_));
  NOR2X1   g1320(.A(new_n1801_), .B(new_n1800_), .Y(new_n1802_));
  NAND2X1  g1321(.A(new_n1802_), .B(\V262(0) ), .Y(new_n1803_));
  NAND2X1  g1322(.A(new_n1803_), .B(new_n577_), .Y(new_n1804_));
  OR4X1    g1323(.A(new_n1804_), .B(new_n1463_), .C(new_n1458_), .D(new_n1048_), .Y(new_n1805_));
  OR4X1    g1324(.A(new_n1805_), .B(new_n1464_), .C(new_n1460_), .D(new_n1459_), .Y(new_n1806_));
  NOR4X1   g1325(.A(new_n1806_), .B(new_n1804_), .C(new_n1457_), .D(new_n1067_), .Y(new_n1807_));
  NAND3X1  g1326(.A(new_n1470_), .B(new_n1428_), .C(new_n1797_), .Y(new_n1808_));
  NOR3X1   g1327(.A(new_n1808_), .B(new_n1807_), .C(new_n1431_), .Y(new_n1809_));
  NOR3X1   g1328(.A(new_n1806_), .B(new_n1455_), .C(\V289(0) ), .Y(new_n1810_));
  NOR4X1   g1329(.A(new_n1810_), .B(new_n1809_), .C(new_n1799_), .D(new_n1076_), .Y(V1669));
  INVX1    g1330(.A(\V205(0) ), .Y(\V1671(0) ));
  OAI21X1  g1331(.A0(new_n1801_), .A1(new_n1800_), .B0(new_n577_), .Y(\V1679(0) ));
  INVX1    g1332(.A(new_n508_), .Y(new_n1814_));
  AND2X1   g1333(.A(new_n1814_), .B(new_n498_), .Y(new_n1815_));
  NOR3X1   g1334(.A(new_n1815_), .B(new_n1018_), .C(new_n1452_), .Y(new_n1816_));
  NOR4X1   g1335(.A(new_n1815_), .B(new_n1556_), .C(new_n1029_), .D(new_n920_), .Y(new_n1817_));
  AOI21X1  g1336(.A0(new_n1817_), .A1(new_n503_), .B0(new_n1816_), .Y(new_n1818_));
  AOI21X1  g1337(.A0(new_n1460_), .A1(\V56(0) ), .B0(new_n1096_), .Y(new_n1819_));
  AND2X1   g1338(.A(new_n1819_), .B(\V100(0) ), .Y(new_n1820_));
  MX2X1    g1339(.A(new_n1563_), .B(new_n1820_), .S0(new_n1818_), .Y(\V1693(0) ));
  AND2X1   g1340(.A(new_n1819_), .B(\V100(5) ), .Y(new_n1822_));
  MX2X1    g1341(.A(new_n1822_), .B(\V165(7) ), .S0(new_n1816_), .Y(\V1709(4) ));
  AND2X1   g1342(.A(new_n1819_), .B(\V100(4) ), .Y(new_n1824_));
  MX2X1    g1343(.A(new_n1824_), .B(\V165(6) ), .S0(new_n1816_), .Y(\V1709(3) ));
  AND2X1   g1344(.A(new_n1819_), .B(\V100(3) ), .Y(new_n1826_));
  MX2X1    g1345(.A(new_n1826_), .B(\V165(5) ), .S0(new_n1816_), .Y(\V1709(2) ));
  AND2X1   g1346(.A(new_n1819_), .B(\V100(2) ), .Y(new_n1828_));
  MX2X1    g1347(.A(new_n1828_), .B(\V165(4) ), .S0(new_n1816_), .Y(\V1709(1) ));
  AND2X1   g1348(.A(new_n1819_), .B(\V100(1) ), .Y(new_n1830_));
  MX2X1    g1349(.A(new_n1830_), .B(\V165(3) ), .S0(new_n1816_), .Y(\V1709(0) ));
  OR2X1    g1350(.A(new_n559_), .B(\V280(0) ), .Y(new_n1832_));
  NOR2X1   g1351(.A(new_n920_), .B(new_n916_), .Y(new_n1833_));
  NAND4X1  g1352(.A(new_n1833_), .B(new_n1832_), .C(new_n1432_), .D(\V240(0) ), .Y(new_n1834_));
  AOI21X1  g1353(.A0(new_n1371_), .A1(new_n583_), .B0(new_n1102_), .Y(new_n1835_));
  OAI22X1  g1354(.A0(new_n1835_), .A1(new_n493_), .B0(new_n1834_), .B1(\V172(0) ), .Y(\V1717(0) ));
  OR4X1    g1355(.A(new_n562_), .B(new_n486_), .C(new_n1409_), .D(new_n1096_), .Y(new_n1837_));
  OR2X1    g1356(.A(new_n1234_), .B(new_n589_), .Y(new_n1838_));
  OAI21X1  g1357(.A0(new_n1838_), .A1(\V1536(0) ), .B0(new_n1837_), .Y(\V1726(0) ));
  NOR4X1   g1358(.A(new_n1798_), .B(new_n1474_), .C(\V802(0) ), .D(\V290(0) ), .Y(V1736));
  NAND4X1  g1359(.A(new_n1551_), .B(new_n503_), .C(\V33(0) ), .D(\V289(0) ), .Y(\V1745(0) ));
  XOR2X1   g1360(.A(\V15(0) ), .B(\V16(0) ), .Y(\V1758(0) ));
  INVX1    g1361(.A(\V101(0) ), .Y(\V1760(0) ));
  AND2X1   g1362(.A(new_n1482_), .B(\V56(0) ), .Y(new_n1844_));
  NOR3X1   g1363(.A(new_n1844_), .B(\V1760(0) ), .C(new_n1096_), .Y(new_n1845_));
  OR2X1    g1364(.A(\V15(0) ), .B(new_n1019_), .Y(new_n1846_));
  AOI21X1  g1365(.A0(new_n1814_), .A1(new_n1551_), .B0(new_n1846_), .Y(new_n1847_));
  OR2X1    g1366(.A(new_n1847_), .B(new_n1845_), .Y(\V1759(0) ));
  MX2X1    g1367(.A(new_n1233_), .B(new_n549_), .S0(new_n529_), .Y(\V1771(1) ));
  INVX1    g1368(.A(\V134(0) ), .Y(new_n1850_));
  MX2X1    g1369(.A(new_n1850_), .B(new_n540_), .S0(new_n529_), .Y(\V1771(0) ));
  INVX1    g1370(.A(\V78(3) ), .Y(new_n1852_));
  INVX1    g1371(.A(\V1213(11) ), .Y(new_n1853_));
  MX2X1    g1372(.A(new_n1853_), .B(new_n1852_), .S0(new_n529_), .Y(\V1781(1) ));
  INVX1    g1373(.A(\V1213(10) ), .Y(new_n1855_));
  MX2X1    g1374(.A(new_n1855_), .B(new_n1041_), .S0(new_n529_), .Y(\V1781(0) ));
  INVX1    g1375(.A(\V37(0) ), .Y(new_n1857_));
  OR2X1    g1376(.A(\V1243(0) ), .B(\V37(0) ), .Y(new_n1858_));
  OAI21X1  g1377(.A0(\V1243(9) ), .A1(new_n1857_), .B0(new_n1858_), .Y(\V1829(9) ));
  MX2X1    g1378(.A(new_n1853_), .B(new_n967_), .S0(\V37(0) ), .Y(\V1829(8) ));
  MX2X1    g1379(.A(new_n1855_), .B(new_n956_), .S0(\V37(0) ), .Y(\V1829(7) ));
  OR2X1    g1380(.A(\V1243(6) ), .B(new_n1857_), .Y(new_n1862_));
  OAI21X1  g1381(.A0(\V1213(9) ), .A1(\V37(0) ), .B0(new_n1862_), .Y(\V1829(6) ));
  OR2X1    g1382(.A(\V1243(5) ), .B(new_n1857_), .Y(new_n1864_));
  OAI21X1  g1383(.A0(\V1213(8) ), .A1(\V37(0) ), .B0(new_n1864_), .Y(\V1829(5) ));
  OR2X1    g1384(.A(\V1243(4) ), .B(new_n1857_), .Y(new_n1866_));
  OAI21X1  g1385(.A0(\V1213(7) ), .A1(\V37(0) ), .B0(new_n1866_), .Y(\V1829(4) ));
  INVX1    g1386(.A(\V1213(6) ), .Y(new_n1868_));
  MX2X1    g1387(.A(new_n1315_), .B(new_n1868_), .S0(new_n1857_), .Y(\V1829(3) ));
  INVX1    g1388(.A(\V1213(5) ), .Y(new_n1870_));
  MX2X1    g1389(.A(new_n1335_), .B(new_n1870_), .S0(new_n1857_), .Y(\V1829(2) ));
  NAND2X1  g1390(.A(new_n1355_), .B(\V37(0) ), .Y(new_n1872_));
  OAI21X1  g1391(.A0(\V1213(4) ), .A1(\V37(0) ), .B0(new_n1872_), .Y(\V1829(1) ));
  OAI21X1  g1392(.A0(\V1213(2) ), .A1(new_n1857_), .B0(new_n1858_), .Y(\V1829(0) ));
  NOR3X1   g1393(.A(new_n1802_), .B(new_n1595_), .C(new_n576_), .Y(new_n1875_));
  OAI22X1  g1394(.A0(new_n1875_), .A1(\V1833(0) ), .B0(new_n1617_), .B1(new_n1611_), .Y(new_n1876_));
  AND2X1   g1395(.A(new_n1876_), .B(\V14(0) ), .Y(V1832));
  INVX1    g1396(.A(\V301(0) ), .Y(\V1863(0) ));
  INVX1    g1397(.A(new_n1021_), .Y(new_n1879_));
  AND2X1   g1398(.A(new_n1485_), .B(\V56(0) ), .Y(new_n1880_));
  OR2X1    g1399(.A(new_n1880_), .B(new_n1741_), .Y(new_n1881_));
  NAND3X1  g1400(.A(new_n1881_), .B(new_n1055_), .C(new_n1879_), .Y(\V1896(0) ));
  OAI22X1  g1401(.A0(new_n1880_), .A1(new_n1732_), .B0(new_n1055_), .B1(new_n606_), .Y(\V1897(0) ));
  INVX1    g1402(.A(new_n1419_), .Y(new_n1884_));
  OAI22X1  g1403(.A0(new_n1880_), .A1(new_n1722_), .B0(new_n1884_), .B1(new_n1551_), .Y(\V1898(0) ));
  OAI22X1  g1404(.A0(new_n1880_), .A1(new_n1713_), .B0(new_n1884_), .B1(new_n1814_), .Y(\V1899(0) ));
  INVX1    g1405(.A(\V15(0) ), .Y(new_n1887_));
  OAI22X1  g1406(.A0(new_n1880_), .A1(new_n1702_), .B0(new_n1887_), .B1(\V16(0) ), .Y(\V1900(0) ));
  OAI21X1  g1407(.A0(new_n1844_), .A1(new_n1685_), .B0(new_n1846_), .Y(\V1901(0) ));
  INVX1    g1408(.A(new_n1708_), .Y(\V1921(4) ));
  INVX1    g1409(.A(new_n1719_), .Y(\V1921(3) ));
  INVX1    g1410(.A(new_n1728_), .Y(\V1921(2) ));
  INVX1    g1411(.A(new_n1747_), .Y(\V1921(0) ));
  INVX1    g1412(.A(new_n1682_), .Y(\V1953(1) ));
  INVX1    g1413(.A(new_n1775_), .Y(\V1953(3) ));
  OR4X1    g1414(.A(\V108(4) ), .B(\V1760(0) ), .C(new_n1887_), .D(\V16(0) ), .Y(new_n1896_));
  AND2X1   g1415(.A(new_n1896_), .B(\V110(0) ), .Y(new_n1897_));
  OAI21X1  g1416(.A0(new_n1681_), .A1(new_n531_), .B0(new_n1897_), .Y(new_n1898_));
  INVX1    g1417(.A(\V110(0) ), .Y(new_n1899_));
  OAI21X1  g1418(.A0(\V1758(0) ), .A1(\V102(0) ), .B0(new_n1899_), .Y(new_n1900_));
  OAI22X1  g1419(.A0(new_n1900_), .A1(new_n1814_), .B0(new_n1898_), .B1(new_n1096_), .Y(\V1968(0) ));
  INVX1    g1420(.A(new_n1236_), .Y(new_n1902_));
  NOR2X1   g1421(.A(new_n1410_), .B(new_n493_), .Y(new_n1903_));
  NOR3X1   g1422(.A(new_n1903_), .B(new_n1902_), .C(\V134(1) ), .Y(new_n1904_));
  NOR3X1   g1423(.A(new_n1903_), .B(new_n1236_), .C(new_n1233_), .Y(new_n1905_));
  OR2X1    g1424(.A(new_n1905_), .B(new_n1904_), .Y(\V1992(1) ));
  XOR2X1   g1425(.A(\V134(0) ), .B(new_n1233_), .Y(new_n1907_));
  NOR3X1   g1426(.A(new_n1907_), .B(new_n1903_), .C(new_n1902_), .Y(new_n1908_));
  NOR3X1   g1427(.A(new_n1903_), .B(new_n1236_), .C(new_n1850_), .Y(new_n1909_));
  OR2X1    g1428(.A(new_n1909_), .B(new_n1908_), .Y(\V1992(0) ));
  NAND4X1  g1429(.A(\V257(1) ), .B(\V257(3) ), .C(\V257(5) ), .D(\V257(7) ), .Y(new_n1911_));
  NOR4X1   g1430(.A(new_n1911_), .B(new_n1129_), .C(new_n1192_), .D(new_n1166_), .Y(new_n1912_));
  XOR2X1   g1431(.A(new_n1912_), .B(\V257(0) ), .Y(V650));
  NAND3X1  g1432(.A(\V257(3) ), .B(\V257(5) ), .C(\V257(7) ), .Y(new_n1914_));
  NOR4X1   g1433(.A(new_n1914_), .B(new_n1129_), .C(new_n1192_), .D(new_n1166_), .Y(new_n1915_));
  XOR2X1   g1434(.A(new_n1915_), .B(\V257(1) ), .Y(V651));
  NOR3X1   g1435(.A(new_n1914_), .B(new_n1129_), .C(new_n1192_), .Y(new_n1917_));
  XOR2X1   g1436(.A(new_n1917_), .B(\V257(2) ), .Y(V652));
  NAND4X1  g1437(.A(\V257(6) ), .B(\V257(4) ), .C(\V257(5) ), .D(\V257(7) ), .Y(new_n1919_));
  XOR2X1   g1438(.A(new_n1919_), .B(new_n1179_), .Y(V653));
  NAND3X1  g1439(.A(\V257(6) ), .B(\V257(5) ), .C(\V257(7) ), .Y(new_n1921_));
  XOR2X1   g1440(.A(new_n1921_), .B(new_n1192_), .Y(V654));
  AND2X1   g1441(.A(\V257(6) ), .B(\V257(7) ), .Y(new_n1923_));
  XOR2X1   g1442(.A(new_n1923_), .B(\V257(5) ), .Y(V655));
  XOR2X1   g1443(.A(\V257(6) ), .B(\V257(7) ), .Y(V656));
  XOR2X1   g1444(.A(new_n1616_), .B(\V268(0) ), .Y(V1370));
  NAND4X1  g1445(.A(\V268(4) ), .B(\V268(2) ), .C(\V268(3) ), .D(\V268(5) ), .Y(new_n1927_));
  XOR2X1   g1446(.A(new_n1927_), .B(new_n1612_), .Y(V1371));
  NAND3X1  g1447(.A(\V268(4) ), .B(\V268(3) ), .C(\V268(5) ), .Y(new_n1929_));
  XOR2X1   g1448(.A(new_n1929_), .B(new_n1613_), .Y(V1372));
  AND2X1   g1449(.A(\V268(4) ), .B(\V268(5) ), .Y(new_n1931_));
  XOR2X1   g1450(.A(new_n1931_), .B(\V268(3) ), .Y(V1373));
  XOR2X1   g1451(.A(\V268(4) ), .B(\V268(5) ), .Y(V1374));
endmodule


